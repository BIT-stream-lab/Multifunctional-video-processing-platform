


module hdmi_1_4b_receiver_core_wrapper#(
    parameter DEVICE         = "EG", //"EF2","EF3","EF4","SF1","EG","PH1A","PH1P","DR1","PH2A"
    parameter EDID_INIT_FILE = "NONE"
)(
    /*
        clock and reset signal
    */
    input wire        I_pixel_clk,
    input wire        I_ddc_clk,
    input wire        I_rst,

    /*
        tmds raw data
    */
    input wire[9:0]   I_ch0_tmds_data,
    input wire[9:0]   I_ch1_tmds_data,
    input wire[9:0]   I_ch2_tmds_data,

    /*
        hdmi ddc channel
    */
    input wire        I_ddc_scl,
    inout wire        IO_ddc_sda,

	/*
		hdmi hpd signal
	*/
	output wire       O_hdmi_hpd,

    /*
        apb bus 
    */
    input wire        I_apb_clk,
    input wire[11:0]  I_apb_paddr,
    input wire        I_apb_psel,
    input wire        I_apb_penable,
    input wire        I_apb_pwrite,
    input wire[31:0]  I_apb_pwdata,
    output wire       O_apb_pready,
    output wire[31:0] O_apb_prdata,
    output wire       O_apb_pslverror,
    output wire       O_apb_int,

    /*
        video output interface by native
    */
    output wire       O_native_vsync,
    output wire       O_native_hsync,
    output wire       O_native_de,
    output wire[23:0] O_native_data,

    /*
        video output interface by stream
    */
    output wire       O_axis_m_user,
    output wire       O_axis_m_valid,
    output wire       O_axis_m_last,
    output wire[23:0] O_axis_m_data,

    /*
        audio output interface by stream
    */
    output wire       O_audio_valid,     
    output wire[23:0] O_audio_right_data,
    output wire[23:0] O_audio_left_data,

    /*
        arc interface by stream
    */
    output wire       O_acr_valid,
    output wire[19:0] O_acr_cts,  
    output wire[19:0] O_acr_n    
);


`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Anlogic"
`pragma protect encrypt_agent_info = "Anlogic Encryption Tool anlogic_2019"
`pragma protect key_keyowner = "Anlogic", key_keyname = "anlogic-rsa-001"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
dYIx2gMN2Jc/3SZxzB/xSB+Qu7bISCIx2XxRotHepzSLCVtK3Qzq4r6R/R/ZZNBM
VMazYhwmAGsWq/pEq7PRAaGoDEqV6qvwRrqi5YPGwdsEUjxqkbx2lZFmuHc8qTy6
b0OGEJDaJRKV07QJgMS0PAlhIYif5Rfxv6YiMCTk/Gs=
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "CDS_RSA_KEY_VER_1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
hrtFEQpCbjMLVHcqh59izKYT/AMPRpviUq//9K8ydDCjuDxYeRP1UBP99vWWaZ/U
3W7GHqtyQdKh3m3I3pNORREASM8JoMHEZ+HZQShXcSufB+Y786rq4n90+A162HGI
l1TAfwFflk9Hh1dV/8vzo+eD1/yOKeXvlGk4qtnWY47uPFxdTMLw/cLedZutdh8w
JPT9L1fEODIQl+lzgBSL08JX+dhijUCY8YjcJKupcXbxtgl1xxCAzG2DmRzcJ5yU
BfJGMS9i2ecmVCxDYahgH+lQSx4Wmr5K4s0vAMUzo9GCznZnQXB8jvUtqo//ny1z
ole59O1gaciN8bnJ8vpoUw==
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
b8dIXEQTmWi1gGA0rsZn6GjEj+BnfmnSsEqWCzKZarIdXVNI3gaOwcsz+jy/q1Y9
pXOniJDWaz63KbJMTXeS9Ghj7kFx8vszGged91yjO2UoMq7DdbSHJ4Dk90OXvztt
hzfmfWam+pYmWfmVXZLYHGeioeLuTQaFjDe2f/FzyWQ=
`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 256)
`pragma protect key_block
faKZy6uEg4EjcEsQW0Nh3GZ7of8YEYk2Vcuq1WkAlPTxJhBCriW/Wq9Bo/j0K7tR
Py44m39jrj8P+3KRHjkEt57qimzHNN2s3J+hbb/6POy32TAIa1L0sKu6HxW24q+Y
0xBqk4x3Pz9gXvpkkCU69NGjVltimsKkYmJlt5F9p0vpeSZZ0RLpmkBGZUf78boZ
6StNLqH+C7ufXQN52Vf3t39KwHHgv59q6wZLtAlvKZr6yW6wGkc7moI7OVV+9QV5
TTRwAblNirqJSCx01stiZ5NyjEt+66MxciIY8B0BcgXJOVGgCEGw2JjGXAaWGhs4
PWsr59wpDV7x2sKEOWAjyg==
`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2"
`pragma protect key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 128)
`pragma protect key_block
ufT6FWfSmQWMO/TRSGLTLnNWEstqbAjeqrXAnGYmtzThvXwbuf+PFAo8nmBqNFfV
FiyKvchhDLWa/4t8SRx5dDMXnak1qawfU6j1+VWhw6xtcK8iS2NMsEM4CtUAuesh
nOVG3394dQfIl+XaP+ueuzmNCG9a3WiPp7pwAOHZr4w=
`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 64, bytes = 200496)
`pragma protect data_block
wJHBlOLmtVzjaXMMj9GCwNjjp/Bl2j8wKRz3wMQtc+84N0dAKgcj/JaOMjzPOHRb
G9FqNp+3Re1+7uMJQMYtJFuXmWbFoPv57MfgbewABvrNGZFV54AOyNq4DYLgkCVK
iHJR9QVJXXXt+GBWdkUpQwuL0xYxjUyfpBMm4qjyCK47J2T40E+sASAUHAXDyF1f
11tz1Yyb4w1zk1h4nf0Fly+dv18iWjtkIzxIrrhBqs7Vn6WGM/qZ4lCvJwUVL7aA
qfexQPgYURuRpuDEJfpS6QncK/5maw+aKhwF1C6Yzr0PqBjkSygSxPfQuNh34ayI
G4dYSpMFEkaHZ1nM1/DtH8Or05qAXtkaDJSTkfCjVTWGg43EGoDCtZoShfqFq4ak
OilkzcLzaujpRzjUv2fRd0U7dbsu3KqDEcQMC6V+0kw8DEb98xtPsuUnvTJxuWmy
47wqXEM+naNqCgAQQO+Ico3u3+Brf2IWPWVTVn1clIvgjxYTQ9WpD3YpL0Fi6dvY
WcyW2WXxNDoYr3/2KJkOVu8nSvr+id2+8suyH98nSaANqdkTPBX6q8Y64+n5B2Mp
vVeKt0F9dOBrTDx8YdjPTeRC5XkfhP/t2glm/JlbwOZbx/zD0YvIwGhtmZBRPq98
Nqxv/6btbqQdzXRhFv6NgYwytxAcEwr17jg4RRL1VUiNgUpaGG/1Mm7+VnbmE9ne
NrlDSLey45DT3V4AK8TYVigrbI7v+AgS6eBwOlVd76rpOekkcW8J8RA4l4kbl8iy
hpqGPS04TiAkU4I7lQ5EKRj2GbGksqaOSvzwSmqSQx1SEdnpt1i+0zhSpC7/NSFH
bPQdlGjicskLq7H13rOu7ClPobZ5sz7lu+ybpM00Qe3lK0INiTRPKXyVZKcYktXZ
z5hMVRodqXsF5tt6jaP72XZ8qWhxBGFb2s5NfqUPCoG9Fve0akM1Z9IcTAEg7Ozk
I2fp+Xeg0V+7ntQsEveRbGSvsx14zXy3NKdOCT/BjcV7mqJsL+wBEaIGLuyHcP/p
UIWwJJMS30kIFegYj2zWc+4lEiYYrfJVMwPjqf/vYONT55UANkIfTFYYWybFw5XC
LgCla3CaAabjdSxr0TNY5O4L0u1U4/IRBXhknkxaOqW7R5FVHBESgcRG57uqtXKL
WiXJUKAqQ/T1a0qxWFpHj0j+bEf4oyqf/bm7w6v8RV6xZl9RhEWsdSSU96g0/sKO
x3lFqZxmUfaGeEScKOSDu+ztDAtgBwttTWNdHxaU/3n559Ws5NLhNspvMYRh+lFL
mv+bBHGzEtUDu6s0VjQUxkVyVlAF2pPRnO+yKBPI34wIMltRv0qOXRAI9vT6Mk2N
Fi0NPbBd6QaDLtcyYEUWer+i/OC4QMGxAyBNzaHWymGfFD+Ki8FYT1753SipVx3x
t4NG8t0qkAUus7qYBAYp9uEIWdRUwq5GkRk7N3hJN2Uy9pshnRLF3kwHDPnAcDHY
x5mjjShHLlPO7+5k7klG8j5xU9KCQug+rucKva6iQ6x9eBnKgZoi4T4R7OOCZXXw
OG019awfnayoATE9CDrvsqjBQNyAMQPfIyj2ZL7So07K038C+XYonDGbL9KaUpDn
zCs7QHdyGey9eHOSun6i6hUqedk+wX6brl7VsJYFZ7q/GAmJL/eUvnFN38Ne7/fx
GaQ2YCpWj0/AkS/Pdecf+ajOjaDGmclhQJXeV2/SMm8x15i32cISf8nSB6njLH7d
7TfjXU+zXKSWe+NaE9APEPMn12NuikgRr3OA6+LETd3Eyp35nDP81BR5RZpq51GR
eWpCV0hF68hxBe4Ziwhem2LWDqxSgw7a6GkU2/MCo2B0UcF8AhlpTImHywAcLXlm
r0FseLAfPaxxoW8k1h3+x+S+8w6lrngfdrO0azyeQBh/L1q+FR9yo0U8tAL/f/ia
wJufcjn6rUw2b0JDDYmxMvODsGWbjEm5t4WkrVkAw3HIGGxbuCzvu3MkO4hZEMRX
OOqNcLJvH0f85QETtPIkeSomsiVSgeHlKIORDGXjfco/5qYiJsfMYZSfGaNTfrTv
c8lnuzn94CjU78N6odnW71MfjLUOj5Zmb06bSQg29RgcAu0INdb86F9F4EXmzwtR
2VH9FaJPG9j/gysA1x+eehRPVGrHAHMt2kWoDNgBG2v6DPcKGx5XGS4iBmbQzBQK
n+FuZVzswtBRSy6tUmhFrpQ/1gBiGqCmV3gwvyo5smMxNwbnGBEnwiKPlTqZ4sMM
XlbAT6fhM+Kn//UC1j86D9TFOYVdiQAJHLaOmKzxjPzSVXfEEKpAEoW13fr3lCzJ
pHwwQShzHnFD/OxcQZUXok4rY4csAN89SFWS5v4xAssp+dS8xuNObw7pXRQ7Gjlf
oQSkho1A1jonm80z2xT3l5j0JtCibapolWz0G/vgSwLJ9Bb87ivqMVXVfurBm0ya
eBvBjzYYM+0Wlc8ee7TDBpqqq71m3vRpUDAU8LNU/gGrg+jW8IqRvhvRfU0yArL/
wwhZQ5wDwuVvJO6imRaesWBL9alQYfruhuEz7jJ1LOVrrPJdLpYBKK5rFOKB1ama
YhKx7B2ze5WQh2nhMMz4a/3XM7x1Q/GWtp2ckB/NX14EgUQko3w4kb0R5uMBkbnz
D7ForEnFMduB4gKuZIYEzbPXVC0m/Z9KViQkmD+A5ZV07GWhTi8jbK9lPAId5CNl
lfxQmT+NF3i9TYUhNA7eEFh3NQs42i3WrwavRvY7WiSPhWwHiW0YKHH5YJTveMlk
k2yiwLNE/7KCVTjPK/TMIFrcM/WkhHFwfbuG2jal+I/Nrd6z+PVz58yfZ5mYlXgt
jCtac8Ns51vmCu7ZhGrh55tfciXo0y6k7Ichlce9hZGof5BGt7hvizX510CQv1/R
FsGGueQr3dP/++pzRazQ9EpIUEoCGxhobC8QufG9WBZ5gtzNM3U7I87I7DZaWQ0E
/CW/U8Vy5yBKqyrhtT051Alq3osWlXMYuXQKwjv/wkIgVXxPvSUyPjV6YYVJXUda
KJZFuPiTje7VuyeHdJ0Jor+YWvZhK4B8Slui17n9NkB5T7IVARS0VMFEj20hbxxl
GiGrv3tnIa/sGkra7XyWrGO7EQYWJVuufh3G+HaggxHddX+tWQYTzKhUAfD6lncC
i9doUiVUvgL+sP//3jbkIVzV1Od5yY5txumcEbb7M0SioaNsivSbE8L4ohtgKX5g
1oy26Zs7krLGhKOjEiSaBTdFfwYHfxJ3K1M+KcZn7c0jwjJ1wk6NswG1zwdE5JQW
+hcPbixZj8APJ1HuH0S/mHnfyN4wPjcEvr+oXIKei1DGwt52O812Q8RoUfveBKC0
0vqGUY5oBYRZpLlsrWicPkRC3m+jgKYBNr+8fSqF/NXIqlM2sDVeWRzpnDgcinqo
xWe5UPUkKSC4XHtKpVxqIOXDErx/4UVeHj67rWIUTrdZqV54i/6xmV9VicwzgLot
rSMiwjKM0sgudP/MLppwPLDIbEVJZYgesjcwH9L47vuHHg7UlDpKkJnDpoAXJ72E
tqHk9FeiU65Rs0w3LmuP2J44AmlUNlwLVAeWEo5iAAEoB7932zBJGXKCWGjurIL2
LNJq9GRZw7NHR884Blu3vHBhLLvcOs9MS7oggZ3th2wq6L8EYsBqbPQgtHPwtJ7s
ssYDirARQoZ1ZrJgqv75YvJ/JQCB8kxcByXpp/VvlC2tUK+uQFcZ6iCMHhKGc8ZV
G3oEo5T28bZQb+b3ckNf5ZwmnxnbdGDGfKZM6Oainh0Ct9vU9ic/aguBoBqLu1UL
ho5XbHFkYfhb8HjIgGZhrJ2V1C60V9/Z5LZhsyhDRv2SUb1+tfyxWVopJZWm0Yps
BOulFsC79icGdtIepLVsGUSCISIaEWCcpMYa2j4iRw0GvxI+1Omaa9ZMkgA7ZWus
LF43Thp30uZmPvjqszkc7HnHWPq80OzFFNbYR21o99MiNdrz7ANt7m3DTX/iZ2XJ
MDpbHsPXit6EC4+oABcwwoAxGn5+LAx8t2m3FmOaU/Bjco2LOthjBtWYtRtz/tZw
limCrv+azFRZUgNLwPErdtGBvDtxOxh+72NRvq0RA1rxygvRnWOmOvBFljQ5x3Qy
5WKloiBc+Cvd31rhRo6ZR2A7xeD+IU1rpNK0TGSpt5UdxSInoKLjWuwbnl9x0UrH
uxTWxeYQQwh1JuXng2+agpOldFDqBooYtoqoTGlfjqDzZDxwPUdBorNmhwalMl1K
hYOrbbY55USItSi8s8IycvAC8ZzRvmYITa4bSqDBn1WLtHXlxRutLz10Wfj7ho0C
omxcOZcrwneWH8LKXlJR6ScY/ponPEVWgsAYBUl4ywcd+ne0owBW23UQN6Ovl4+1
mmUjy1Ypu4+RsQWdK1Tjf2l2H2uDCULNxhVr0UMyyJaIIdBx61D/nxWQ+Wy2xFaY
+ekdAMfpeHdZf1w5yuGLSbOrE8ltqb9t0VxibvD57VKi/swHMtPJRw0qBcNr3k7G
dME9EP2FWghcg8OG+WQnxUFZHhDI4+KNQdkollR0xVJ/TSt9kYFZQNvZN9kQsrtC
xullVOnsTj21c7G2cyuTd7ueZwWVpdoXHGOsrdgF6UwNh8OtNzvY74Y4Vnt73piU
laL0h2wMgkxr52uZlGfQnpbh5C/FbofgR8Mmq4nXacRrwX/hL9y8sMNcb+PaQMca
34LXQ/I5j8EkQXoCtZfY1CE+8iPuAmo9XP8vJ2fmizW+3a9zIvTQdNikXYEheuff
5v8lWYlt8nPBNtsnJtj4JhCxFlGQcA2ppbfiaaHjQJ1aNfkuX+FsDLIiQjtXR4o1
O5z3V10HYPtJ9IWs1tScU63LH+Xie+Y0RkfrSe5YU3P1/xkLIBvZxJ79Hsku+5cz
MQEVgSwR+x/fIIwYOSJez74POTujYpao0klff5IuusO9TLDDXCaeSGOCVKpMprS/
2opaf+t2SslOHn2M9YEtcRfOnfQdiXHn3TaMMdxxw0IlNpD5h/6wzVyeHxdp6Ide
tJjSLZwlxxI/KfYI8ExydqnsScjIdYebfCVysvephReQFSjAunr4MjZMzt/O30ba
U0s2Jt0pS7MfLORfv8Wf10BcyEGiZV0KpN3CBgaaIUm1Yr54sd37DVajjEovKmDl
grOCKuOt4nwDJTDJuTrnK5ki2BImFix6bMZHUzImFdHgX1UFDHOzmVOxuB+2Zy+V
B5l/wpCUTr7CwsAMaakNu4yXFFSnZsNsvEUwL/490GOQnhj5A3TAnA6wXCw4KMnA
p0LNgkqAnRUj3C4DGciaPac1zhF10PiC9WyxyotXCFa2cPaxXYDSCGCcPWHJpitm
J2VHie1iR3Si4gpp61NmycLiS0xbvRTf394hBkcFKbx5kHbH0X8ZnmuVESYPjCxF
Z4OfRb05+GyTfLrqk5fhEbebe4M0PhzIPQBcPLyCx/l4BKd2jOWzEg8ElTb+qNRM
twSzQhoO2eD6gQN9APXYK91vHlawrJJ59iP9feumBDK04M/p7CFYmt4ICHucCRii
LhsJy9t6Z9rNlbQuNbgQD8hSImNLL5uvFG8Q2X8OQd87wP399XyjUdxdfy8gXczB
SuhfqlPn/EG/0jw1oV9sK8YljCIlCzkWPBEKAKaRi+Jw8nuROH3jfxoWHh6ZE0v/
dZHIHE1vdLvEVCzoxFWsIiVMwaeLetZGpDU8eZo6QKAV8/ukCcA437jQTx/ywPym
v3aZ+84nbHhAxUR0iYcabEzwpHNvJOYcA+k/OADQ7n+qzEZ2LJ5bwxpo5QHA9BZA
cuogcpEVMLwaJbSs37eKJ27oK15+c2pYAH6sqFqftbVqwl2I9/dGU1Clzz26V1TU
srp/rYjmVQH/ko1Qk7uh1QNTJK766RdjoCdNvpY5j7jCCqrVZHDvpeGTSgNleLOU
dYvW+OXk9pW22c7HoZORyZm6Ex4NDZ09hajRDxWCOv+nka3y7b5OlYQlYnSnq053
5fprzDhpAaUzup9yU1Ilmv7x2xeJ0D5qimMElgtFPVBnqrjnxPn+apzpqCZU9pSR
QDDzZ8iwZHlp7wfnUfG8OdmGUAGW2/sX2QR46chQ/4Yf60DXRucSu42pHEjr0fQg
qWuDKvKtIl3hPxuo4xJVWKz9stG5Q/h/dTmEcLIdPSOjgJ0WOoT2GnAdE+LnhENo
ZYaKZhmeur/d2UrTwxdb4bX7ipinlt/GWqj8vhnqth8CeTzRD6Url6g/pmcM9Svz
JhnUGSs2lwWvQdH38R0Ne1x4iqgaGe1mRsno1vrHn01Q/2uFrjTTS0Dirh4gTzop
0BOAPbREBWmDBRTUq1PkPpWpuwV0VAT/u6f3fkAnfjVF8PtfP3qZCWyM27SVCXOO
h3erO2iIeM4xbJRbZR/agQMY2EMaplbuxv1ZD6FhIx1x0Jkv7SJynGiTARH/dulO
oGGkz6QZ9Y5cNmxJAu5JwKASGlJedHBvcW7X4HiJbrO8HIJLGaVq7fR+e/TTPG7a
Z7toaOs1ed5NbZRFmOzQ6ooXLalm9AVKQaM9y73ZQ/bTiHrZmfXs+BDErnDTJ/yJ
tOvhRkK05gCvWLot+9SpCOZU4+tyAUu15tXEPT1jf/CX3crkBjXkIfaw1hl26s+Y
wUnWl+1HffAtV3YtA98uc6dC3ZP4Jz3/Gry66pvLzUtWKSoyyNJmsjv+ljrz/kuQ
3TnV7KVRGOIGBDV+pF2CSCU8Yl+AHzeJItERwAhjmhqPuZi6HEhPP9gRkYIezzKC
uP8SBKN15qBaqu+N+2Aejhp0ZcS4tI+nfIBx9yq8xY9r+YssowDrm+55pf/ob3g0
V4OF0L0ZiMx1L1SauSSpjp5BfnAqFKW7IymoAxKLZ8LhYtO4gmTq4KvItvzswTwG
dGeRW4VC4eE53mJLb53p8hli1qibKUP91ewJPQzwAgqHzHny5k7d2Onvgv4Hpsbs
tDdM4VNms09nZisJUEui4wf8G4lRvlMPFT6xnvbyVyQ5vyV7esMm3fiK6moFHNhE
Mvjc0KMY9eb4NDRpQBc66oZHN3Mz1D5vxShkqqzbuJgv+qxXHE2aGHbOHErlgZq4
3J7LxE4uv01FGt9jNFKzP8L0L5hqXca1GhTH2gLcO5DRGBgMHAvxs2n04qvFT9+W
pTj3nR+M3qeMU9sPIKiSyJj1oVA9DwO3V/ZxnI2z/DAG9UVOIm+AiM7oioxPsYoR
aSh7UIpyXlU3sMzo+qvm+Go4IROrxw2fb4WbcHh3c5CQxrFWiGW9jADiRMBARciw
3V5I/Cj57riCQPWh5d0yGXT7m4I7psPYCreFJbdr/w+UfbOwgOSrGpQTd3uCa6s4
BSOfp/zgKGdafJ5AvGsCkMhaoly/OGmc36zA2paKkWBOG3wBwy784uWNCLBGVTLy
hXj6h6n7Uq4JyiC8InAQd1nCayeQpmzZ+V322XQU5pQb3w8Z42WJgRoRN77OBUPQ
vTutAPlh9vzvdiP5+XvC++RcJMlQrw+DPEp6IreyEXNeGT9Pt7JURfdgmbqTvC/k
Lqz50ccDcwtzH7Gs7FS1k2BUaJi+SAu29YfwrROJfN6j7ralY4b03+TvpgP0oBXi
mP10mfXiiDGH7dDgzcRl1TrDXom74Ol1b0kPEI3l86+h/D3IEuDMp1wxZMK30d8s
ysm8Ej+muTMAHZxg0p1kt/UNtYXCA6YB6JieX8J2BZZCbc/hnWU8gIAYqDgi1BCN
ZmTf9yIlUFRbwtQtnUW1v4erAnC6/rSisyKBut1629LaxWgLISDpofn7K5URVi4D
5N17F0wXX9Y//2EBMmQJWP1/efvSBPCl/hJ4w4F2F4GgkKMAgOQFc22ujj8gvpkI
7u9liIBtbCUDVkZJzI5ExaJ2R+hE01d9ZV6B8mCLEGz1l8VTMGE7Tl0apkFqlrQs
HvALocyBGIDS2TJXcPxMhnJf6DIscdOFxvSR+SJnJe8tWz+xGRVgiiI+uhoca846
aw3wC8wRtHzmobzgDijvXIwh2G/kyJaw8IPH6iwlHCsNiJSNYQz+q6fVlo2tvFG0
Q/iF5G7lBzJEnx1xDqiD+nSU93eDr0cay1e56u63B4M9mPRimq+dhoFMvXvXgRbn
eRnDXnFxnovP5TxkChlsSo8UxE8bqbs0oPnkm49ID+JSuxAGng6KBDhN03u1k0hs
nMLynyN0BN9GAmsvEIyoosonNI1Wg6gWXLtVT2dGyJJ9zHZO9MJ71IO+54Zjqq6g
gs1pm+WxYQWU8n3qMYk8BRyNERTKY/ucHdHA1pQOWsqGuV0HKvQn+6Nm+3A/FNJT
DCOv8v9CBkidDhItGI/79KAgZ6BA0mMf90o9B3uecyDqx/plmaCr2UxHmZpyAKZe
G2EUKCvlAMEMGMwIe4VgENqzJ9PSVHWuiVSrpleudeVXASXDcuEVKyId/HSJArc2
7AGqa+MgkB5AD6cB7bAsXg1fO9KIH26gtQKJ/grYY1IXGHL8UqyQORyCp/6VJD/x
vQUo7e2CWkh6Wd0VksvyqZHU9zuXEPdv9bM5+LxxkInaMZP8BCiBHOwTpQ8a2Fgw
YlVFX+EjrjxbEkouItPVAy5BnHv84I8ajhD657PMlDC16mdfLz+6PcnmPFRexIG2
0/esGITL2CKCqRRYVWQcovpoTJkB7FHiZS1TN2M2+KcAZeoDLT1UwbJwvXv4iGyN
lJwFgwr3gRuq06HFg0I3pSu8fKEtz5wjnFH5+nmst1MYmhmdheLXi6KTwR6Y4Oju
7bnXHzF+M5QbS/CcisUNdrzQ6t0iaWrAlGWiJbm7vTXZjZBAnv0Ufx7oa5Ww+bnv
zN72mNxridvE2WDGkOMg/x6eGYJ3AB4rjdH8j+JZ3yHtoJkEMWm/jrhu/1Iw8eCr
qwGcAwYOXPK3AnwM3J4H8xgtSWPpzO+eOo+XwUwJzdqfEk/pw8L8MXXgDC2DEOqw
vLwTTwD/q8Xw+6XtNVsJBWE0bpZV5GbfdQuiUB/KoIxs7K6/eH/0MkdpRUI/UAJZ
8+2eQrOI+raFHIC0D0/5MPTAlxntHDI9D84c+T3y/vPjcGQhEizidW3s4xJzxSss
YlEXHdJQUkfDj2Lk5W26egB4W6wUERJlqqv3TK+Cb6wBps080iVaLRu2JfoEXpEj
+wY5gw7dm2zngrHJybPj49diVwY8QzUoal+v47Nx35Ngeex7M2Cx+gho0mk4+cIF
IZkSzSkjIzdanmnoKQ3sP8UaeJK6eFxFAubblf4QhxCWvD1wTuAVPHmVXgRWQSFy
y1i4AqF6X5lngr55ylIsBDp2PdCOTQWbRDiDjUICyyYtv7Hu0H9UTEprfBlFp8ou
8yXlMc5Hsgp6kRj+T280h8bTJkr3i4/Ruj2/S7VtZxq8yD9YxPih/IZsDphEGuIb
AF5t2p+GoMzNvJRJPUsXo45WgxvxfGIyJYrRBWElaZnfExJfqKXgZAvFn+DM6AT0
2tjm42ssfvDeb4fQQO3rnR06jNqcEyHVuKqpITCbWj7ZzhLwRzg+Fhzse8kotRpG
/6BWPYNRVKYeNHQdOWE6YPOJqC9mJduMeJukfHgwmNWTD6ZylNIVslb1fythrQNm
jd9OMqoxG5ZzK2MEZeF7ljSopV4sgD6r9fQugfN/e+rFvYYWPnyGcSH0f21fOEJC
fdAC8RaNGaGXWTgOiadgSj/3Q3XkeebDzS9Rthoe3bqBNDwadV1nsZbd3TgAHAVr
7B9rOtclzYmTgWD3h4Yj5Z/QZq+hQ2dA0GMitKZ1bVTSZrn64AWeZDuhjOvHJbF0
wsgFrwry60I5qDBPcG5/YIaAOwj6HBUqb1j6fFVUiU9NkTBlaTsl9BFI8743UkvA
6FRhi2WO/+ifF4xDN2ivot9YTqfDDOn7UDoB6S+uvWYdZkMWTMRLJ+Hwbzeo58dR
aNEwePrnxF1ZkmbejFdwEJrgYprR8Y6csY6jhxqEbktelf75uPd0RPThRQ3Uok82
v3RqGvZdsOXwvdgD6lWvr06XcYonrljGdNn+eQ/F6z8BfRls+OqiIrtBXbUByYvL
klQHZtNxt6vjwWJKgjv8+N1jFZi6mn27nYmcw7x9PgTJQEonaYbYBUa8Kgw5TeUh
/HlY29An9QwL39p58CY6E4VUBwjQCqe8pOzUGQcejSmuIgeuyFALz9sKuHPgyVnX
n+5egnUup24/cIs0LWmCr8yfb0Iu5/lrNCHvXjrMbtZnMRuv+sgoLF1XKTx4tsKw
Rn3Zd35TKyOSYOCA4ieZQwKmzAq9S8chjx1FqergzeCV4CxTHTt+359FD3nI128P
Z0wUjv3OF/qnKo2KVaHQpOj+OlXrMkDhVzCMx4Tl/QNgEXcbZoIoXCL1g2WYwP2B
LI4aos3cMIgEp27K9uy5NpkCA+U4xz0RM+iAesJe3lWKI21wFKn2yc0jrqV/0kGq
aNNvJt/VTdvPrP0U2WpcbSCC+/bqABwss5i0np8QUs0lmc9UWldfnGsrjVYeHA6C
IiWiMDsSd047KHTlu63Ljk2Jx9t/g4dSWhCNcZYhsZPF2Ta5QQxJNvG4NdWkn9BP
WjcdwKgh/8bbQMt+pullcxaRbk5CxTqFSAE7tbfGtOAiIBS8xq1NnTPPZr/PwcgV
lLHGiF857wfA/eR8keRuH+3BDG0JA2hN9CInFaK5Dm5vaVNxefBVTytMBA/e0fXh
0TC50Qw4g3ayX8qHcHzXdMS1jREF74YDe1JujvWgg4ZCZRcFNEo+Dnj3oYSUlRJt
WeuCK2Laa84c10cyfnzl7LmXZd+AvFsDCH3uXTrkBuDPd2XMtT2wSWQ7t7MUdjt1
4NCFY8kt6y1/7GzmAblxXboSx85/HqGThp927+UqC7OT6aXYhTk2+i08xDQq5/UW
K0ywltww4XcucGVIGm6yNBGxKtkCc6Fy7VTo7ezgDkFnQQT8K99pf2QPdjubj11g
Ba9vCM+F9xmlJQc1IGSzQtOrTuT20LeUxFakl2W50mmYRInrJs3EvXnMKCrVyw1q
hJQ3/+IHdTn6Cp3Wa9ZwnZT26FT8jfRUe2GEMv1D79jV1tvVvDpmZZUQX/yvr58k
UMb2awfsOx1Y4XHK/xzNNEjEM1YEa433Rz8oP7/2+JFZaFKNh03Fa0Me4xeSwBI+
CXWmNgoEBDMPCWbgdIlkntAyW7vPVG1xU9NTOG3D+xMvZnS5LqjzM4xW+71m39io
TSP1LxdBOmDOTS8stHEdCYIDljJ4QcaJ845OvIXuYmmvobJiwXLO+STe5S6oxDoS
S5HzfXzQhssRt7OGgiqkhmQtEOogUPN687FXghuTDqXd5GjrI750dRlnmTbg1etx
+p/7x/4X8tbHpM9vMt/OSD700cO4a+Ushedd8Fk1qQ2YkC0qkRwwELCJibmzuI1K
I70ZDO7TlXojwLEEW9+T6uv4Uka+p/qCc5QX+0Ehjw9+aqSf9IsqvbxU07jPHb7H
aAF+5DilISMzMSzaR2TkK8kDbyxjZxsrsArD9W/4H/Az65Xoemvx2N4v24MSw5R2
BKSXpaFi7nxqTbkUbtUlqGecLPBHbb++G7cwDFVVcsH7dcSzwG/sMNnUixU9N4fZ
KLVseUI6/8dhYD7mfVlnp9DwBIvH30w7SkH0QOt+QW6Uq+00CxNorfsbe6LF2eV6
oERUMtNX8t632nR1DOOcQ5/lAkjQj+IBwr/uBRKigk4oZ+LM+5pLiANVduUvH2o1
JCxvzy8MFlmM3fxFpgd7eRGQ705sYCMDfchaovM8zqa0CdcUglqV6z6kNJEmbF6k
CZRofGpw+g+EhRsYvHpDRDKAuin2d5WJspK78dzvdcWpwgFBdQUDr3qPYsqSdF9o
XRVNI4RsXDrLqPTCa4HXeWcfofJBASAez1BRm6aXCdJj9ejJwZSssUDcQKb21UDa
/xnWoF9KgzDmAYigm7k5kIXa2PebRdf+R6rkQ4aP1EHxSZceGw8Ru0B0vdMNqDqq
BRSOrg/Z/ww7MXs4kYJyxQvojoAuuenGcsNvWeN2J60/a7VT5SSfvcy+k/edxngh
Tq7fhO8u4HaUWB1X6Xat1b1CYMxMqoiZmoXy8uGXWoIP9iHAZzu45eLKderBVmcZ
4F03pKHiS8+MQNT7JXjWOh5c6Dr1aeMzL8bdNWnMbpMvHc8gHVyhRbvWjzLPlz8h
UuPTDJVnydKOaisua7htaHDawciTBkvynxVR18yuD3nBA+ePV/R2W1WNJWvI9t1w
B/PotJMF5YXgNkAqzart8L4D0uvBohWBmpTK7HTiM/1sKq9fROv5QuoAoaFY3RTC
zcT2namDWZwhP28Pb6oMUMbJQ3fSktl8iNjjwfoWsij051It1s74kbPjKgAVe3oI
wb421JxnpKn5LgS8B+WABDo7s0n/qeutqjta4Jf8aBAYTvKzk324wGk+u73ZBpie
ZlICLWkVkt+V5HXRUKnPklE0ugmG/BVlMLagVv7TzJc81qYjMlTsieCQTC94Z3Ck
Ma5jzZz5cwH9ieqFgFSkbfqvBd/jPDYAOdSl4CwUGIZXlYpQtj9cQ0niCohSDHwk
jjm0oEiISm7PCzC6Pe7W2gfhspsigGJRnmFb8Qm2es0eDwwi3cIkxiQvVqc8A03R
gd0EyqYCDh5Al6KoWcDM6Z3jc5RsGN5AMHwkPI9HbpLGYOq+LOjQCZIsAVxQeQze
8vV/s+gIdwn6TK+HVkdDX6iFRQeuHT3wy2NYqByMVvZn3VjWhms9hV4Ug4YXfMj1
LCM4EYZSBKhybAG4AodZGDtPYd3n48+H9EN25cxApewfLcSAjZ1427cOjJGOuBT2
xDiKX0HdmWXYbGcusiW7FVgfpu5hJ6PIwo9W8uRr/9nBWDhmkmNoVg8X/yCYbTdI
THrJeFfMjIUK/mC5fmu3IKp2Wvl2YtLY/lGsG6iBv9xum2dxGwn2Z+kMjeTyi0El
8vtpTr1AFRXWRCF2YBep8i35vvthI8NfB0hPivkd8WAsCsqAhF+qNcllkMz/gh71
57Z3xCWU98+oQBk5yLustslW5Eka83O5auUsJlyEQ7ExVrDMJsxjv14QBdLvw3TU
fjXiC+LN2tTiANVzknSUsp89E687Jv+V7a8QkKsATC89Zx4Kpwbf4PZd+bmvdjzD
CUzjkLy9aAbWKVDB6HLBS3Ln5z9tKM8eNIhXYEWH7a72N9f3scf7EKK/gmPfvXo+
XpROL5S1eA48aGeQhxDwSQCYMoiiCiM1Vg1ewXXnwsU7Ih3Nmg2oJVHhDgvjRGDe
YhfWGggIXL4X9OVmbY0a0DyVivq2j3+z4pHawg9I82/tP0ZZoMtSmomIW9i6DF/G
3Pj+v5jsiXLTzsq8ySrlxr66Nev93Wur6X2AUICiWNuJZv5gZ2beQzqCs3EuZWkF
sGm9cBB0IBCa6uWd5gxesEpiC3Bp7wLUoYv63wzWirbpYsX2y2uXzDrV31kUWHQr
4tBKX/UrIgju8MGBN+RH2CCz43X5pwoelTyGXZ34A+NaQeugunle+AmuCBP+ONV9
3F9ZJhFzqhNauDUIuLkH96kpz8RHkBRRNC11yKXQXTkxEMXN6QFh2yxnlfZsb7VG
/Tp3YMK/I6TaJMAoNi7Gk5DQvkjSH+8elfEIhT2YdIpGJeFT7wbMgG85fQBWUzGa
vEl1HTtvt72V6nAUXY5jrrgWM2dlVTfVj2BE5kpYC6YnSb/FkK4U5uaddSX7RBF3
sEhhb0jzfEninh3yyihgaRZtswBXQgzHEgSYLV5iP/YvQSXMo5jqO/F0xe3mRrJR
ZCdlVwoAtHND/s/CjQcPugTQZM4nx9t+rIZc4oOYDg1vODP0Izn+r+eJjnPTAIrc
Iuwc6Af73Xkqwi4DtiR6InRG4ixeSPvAjoLvPmp6HiAWB6A/2CRMK94TJK4w5fym
zd7WU0Ilb6F+FR8WSqR/kWlS9mAUhlfTGVzt4eA+xnCOq/h27qcJjceWDzGo/Aef
EU6W3+1D0feLhrsBdQ6zOThyrOmu69tscA40DjMvMBzpVvu3h7SYc92u72TXE6J4
TMkreBbqBdJt1mDOe/ouJ+mUBBjdVgA3+7xjxa7amoUzGTppOS6/tQ30iwbaR4OU
t9y7vnCzVZCdpax+Dnh2mui6QVzGOMg8fgWkEmi6r5klbydy//47fCXsd45cMg3i
2/p8esVwTB2Y+jyKqqQ/Vs5pZ7/fNFPCgrtmDPbimHqZEOtEnsPiC84rpFP8RIjj
75eSgWgTdsKDF0KhWm2IUGZQjQqDAGnJow5EDt7MidxY9trSc9fQmpJiFzcv67WD
0rO0vS6f+fYn5USBRF/DZ3/55hATlyEusBEDn9ZsaCIHQBq0epmVzAXcFnEFLiln
oUTcJBP63Kta4f4JDyKzSAs8myz89zDUb0APHOe7EkTId2OHTwQlfXts2Qu+s8Gv
emgun52Q2uSqJBGxGUMiTcnRHVmesVRtZOrkHxznV/NzfuOIRXPm0syMpJiKDet6
6qX9s2t3HXfOoLE6/ABLQ6CqSF1Fsie6TI+IL/tYvSNcJY8DP7DrbNS2FV9TUtyD
Vf5NLEwC5xIqBJsVaUIUThECXTpQ5gs+N58iKMnhUvodHeH1qM3N9ygKf8vEGo5q
U+1OM1II3McogEEjwhONNGW1HuUpHhRkCSZNoTfU0/kigghk2wNUwJqTpcnHPO3g
uGPXTdAyAuGJuqGiftwhjjSxKeno0yphWX4K6k//B4dv/q6M5cZvJ9HJk0ad/E+S
o8hE8fqAehK5hRe1vbrUbpxkRo4ZzJiQ5qVmfdw/+kpX4QXljDrOubm3OAmwvi3o
4JAksJ1/sTU4hP6iGKdheZwV2YaHkEBkCfFjDqrPPXPssLZ8v7t+UmMQyHyk+Sib
ujpXMUEnHuHzKB3EKC0UF28Sjb1qi1m1EAay+nB82cPnzKUbtjuFJ0acLqyO0/v5
dqssm0kDv0mduG2vnJi/xuovePRbo0SznLjM/cqDErlZPR7hjL6h9yHQP0BFsrVU
WJhsU5NBXWB3HTqZ2dxKSaprACnJoQghplsTrrRI85MLmRFieD1fOwAZjW4PSiwe
rf5XcapXJ7SSxz7OLu3xR6OD3sA+jufybclpBEFn2pR2neMDuHF7BQ64Dc+r/u1d
9UNiXUQADKkDXLyJjZ5sYVrkOxiZAOCtPuaOmmT56StZMjMivrflBQOjWNZbfyrt
8oPxIMxE6S0dbF+9Hi6WKw7oL7PzeSSlIgzF7AgmOrK268Cl87uYexcUwCy12WBk
Ze0KwiHXvpxMcR59lkb3p41Ry3EOapYVdKcu5ZJzhWOBKtwivtQPxu0lyTsAQsJ3
WS9HdtxM+kAg+dCs/WvLNG0aB/W3sol0xxNxbieLXn2j0gD9lIJFC94QptEWNhJy
BgAa/qMh/P0hWpaMkPVQtIDn38r6SvpiXxEJfD+zewVCcxF7RL3QEpzD/OIv8j6E
Il0KsnPDj0n889K74MhsCjsY4WxkO9GQWkECgku36qATW1eMTyzO6JxsbYSAL7JR
VP8/Ot1Hj+6I36xyk6zsUbcULseh7Whk6f+2CMdRj+oXpioaKfV+wkDUH8Cm6dJX
z8VELcaullnWvlsP33B6tfR5opvgM/sabkD4OWvxrbXQ4oXb/ZKMCIfOAU2dLVlJ
EvAZzCrOIcCGWUeqCUlpO60SUzX9VazLen3HTa/9XDS1QjdZWT8O7TjaPIH9uErL
jKV4Mji3eUBx7M5BmG6u1XDxqIlqrQz6s4Qzsksb/7u2rgEvyJOKB1QcNvKjtcjI
wNJg3r2KhGzZiI25MbCsnJE21hM2MssWXFB+LXunbm0fIZUGSUs6NRWHDwgcZxFE
TV7i9tSM1X5LVuw4BNM5r0oBa+cfHp62ht5rzIbumjeqNDEWXwXX0669dxgbSkfl
hRHfU7n99GU4HDns9Mea5dVbJMEMPUiBnH+lcoHkKKxhK+fQVg5/Ox2jajMB+pwl
xabGms+qeB6wu7pbGiYYFPmW1li9etLj1SvNCEO/QM8qk+7pwLVYYTM67yw9TsoI
XBJ/BI3jS/cuq1McUOs/Ypq4VPVWkKpe5Ppep/upSGSG7F/YsnhWMu7x+E2x+0xt
5sEK3gEQIzKOByVlYHDcIoAucPW9JxHJPJqUQMtRofGVIXN3F7dp//otwIj5XJg5
oOhFd/Kafrjfic4Jqdf75eEcINWe78RmASNYJEDrrvaJ5QbiXnFF4VeTmyd3gHsO
RV+Q+gxCrATGomOuwxjrNlSLjN9ruVGVQZkhzVvRUDHC8+Rsv6l1uAi3KMOzmsDD
DaBNaSo3uFcWgs2+UAKvq3bm34Y+uxmOkwOG5PH35tvx0xNEjTeIubecwe5i21jV
r4V5K+q7BFTDeyhDAZoT+BESZaZ8BesDldmMWkxZgF9xWG0lQO9Md48nFmMaPpNi
76wRAaM0K6/Gm422lXWkT8Wo/BxbVCnZcck1QUJi6g4L8xT4Z6er4x46xafLpABF
ppaZvtNRVVWykUJPQidIvXG82hZAwxl0NUy4dggbG/QyM7fySZ1LROVdxZd3YgSf
429AKpNPQRTVPMn+aXtYhpjamr59HIbhqk4oLg0SYXrcvQdPwnCrV48MyfI2x/Qz
ONFSMcYFQsUtFeSYpEFJ7QMHNaoqIQl1+ElvBofD/+8KxL6JvbApgjgF89Ntdlid
dYTOom0Tijjt6ku+Vog8SNOAAmgKdDjHZS6sqJNg7fxXGfIICoCEk3nQHgf8sCZ5
kOd9D7AzEzXCTcoPwQeQyNPD0/x1OHV5pBtvxZOCfYKnVp0MNYIZjTtbd8fd5Ci+
F4RbilCT+F3TUtPu59Df3LMOW3CsW003xqckZZSW7c2UB86xjQGqIoEjlueflnHt
9WME8QTPYSp4G5OX9qQ3z3Tc9N9RtLpucte60t0xg3NNuuRfz1TYJrxlanNbpI/w
F89n+z6MVM85DeNeX5kQ1pxi0MfGaV37CCcHqM52pafoA8zrSw7o67OVAv2df+ye
V8tZsHbysLrC0Lu8KKhZrvasPrlxxPmIARXcojMUAUKmCsg7CXj2xB3UqfCjKZUz
KejyWZz6ijrqIQyF7MZbVGunaBets83i91lViaxCcIKK1Rni7wH3OeKedaOHOsk4
sCGEaNzPtEb7/6EnVAfcBJsSMEEvlz9ebO//PmOEEe4HW6gLuIy1Ks3gZqutSPgx
HfHloSG84q5ETVD+eLpZBCYTcpBbPL4dMCx7e236Xz08dye8FYINn8gLVT4Fv4Yv
FNCD47d8ae6dDz/L+vexmhVGWNm3K51jZ82lX9nmIP2wMB5fVI6BzExhl0TRtRfz
q/6vs3U5Q6FhRBs/lluw4abb8AgMbP6imTRw5cmJvN6zCJWcTIULKirAOOgdS6M5
GVyXvp+VK0pYq22c3k9+Jx+xt9O4g31c6Qz5S4951Jykkqdrzso7SR9+lob8zSTP
y/cxzXBjg+/ont/j5EyN66p4xlUqVl6irMMyWdhp9Ki5nSl1m/rEK5oWeORe33Lb
+B3YHTYCVlaog0FyO+F/0q6ORNfjOTOWFyUtRt5Ikzv/HimjWUjfepXGlEw2oxXh
YCfjmqKaEIjKpjO90Nmvg6M4nw9V09EiCR5FlmlGQY9NnxVQnnCG//C7lYD6m8sP
nI2YDO1n9GYVZ5w/S6wJHXl1PEFCFHqmTFRJmPkNBhuPA0p2r3773Ko09wVdzOwW
SbJSeYTOjRD75m2qofeXd/S5yKEwFX0lgm6vgP4Sebkm7oGv1avmnth8Mr34UCxp
UF1bF4E/ZF2H8nhg664pitDyl2rdhNxJzJtKLlFjBW5M4ohTS0+Gf34N8rU34P8R
SatXpapWgh9eCFe2sNI9Yxa0mS9sHv5J4m1TnOZs6hX68XMzEu7MUETfhC8GD47J
TUGaooNwagIS80bnz37O6zRoaV2tkIXQhCqk1DI6SJj/r17JY54amZVaUCD05QpN
ZA+4aef3TuaGmHabfNsy0dwbQVy36vPNW4cN96OuRztHOeEInQRlM2Wv6X2sQ1VQ
JCdwH/PH6Y0MEW2UP3cBTatnnmKojG+OGV/+pBdbaAQjnkQLKl9wucY4TnJtx5nf
K8LYkGF656s89FwMRmxPIFcVC7ZMKOeaaIrKSK8gpRli91ZLPHKRe7inp0+SEPpS
kgtiuXMMPGdnDFpbwXOv0zIw9kDa9t9CUQEiCpdpgsJhTuprp7dfAC7iZ+r97qok
V3ncURdv+BzwIAPaYyA+yTQE6ibftq00Hy2arSWciUnfHBkDv/pfKKJtq8Ys+GuI
apu5yj3db0lg3OvE2HVMqt1KF6TMfKTTEnb1duN60wlzstWCvnyBXPLA2xCB6jaK
eL0YKf47u85bbKGS4ktg+v0bCy7QSAzsAyUqBSAyfjwVetCrNtUpe03ZOXioE6gk
VRZkPXoWB7WnuELEnkJJq8nYwyyvjID9uOWRnZ1PL+7SyOPzHRtyVScVqGdSuXgq
9sJKsdRfFDALQAmhbjpdpMuqBVUn+Ea4FWnpndzgJZjI1a8wXVJfEv5iBidqjOzz
sUR/ImK4+qa4b8YCeHvyhT7R0wajYjIX5w/3grsWtS7KHtVqlc8lp8zNmd5kYqVu
gsDsME7dVV3cpebpQ0C8VhRsFdnIHZq9mqD+dKm6RLbxdETPaBHMenxm+gayYZA4
Um4y9noBvYwqFX1iSraBZq3zHFTTjU2MHsWDLC6B0/+XW4VwCshUh24QPMHvKDYQ
+nXz8rXYRAM/auuulltAtT6hYwanuNdZSGJppZ8TjzueDwFqsAizalXLZUcqMuAp
W0tTAsZXlF3MQrPXSfCUUX4XL+TnG/w2yKFkf1yFjUjGL1ccx/hJMq5ErwslhPyu
xuBy/JYtFbe28fe1YOx9NCt8Yb4SthpNZERZTDqaW41QqdB131UZWRSt6F9Oo+vr
1HLmqBjWK19+5N/5AZMn4ZuIM7mYRwePO2VORypb+aSGDgtROWVVMfJCDDhqcfec
jwPT8yZKT5EQs9q90au9Hzm5MSDI9DvgAEVjzjL1jDyioyjjxyjllzZCgFxRJi0w
o6r0joBs2zz6wg59TL8EoOAEK/oGG7+ql8T8kne1ANTTeXD6R2pwkQqlRpOxwIIA
dLNgmEROajG9WcUNbnCjJOGAcshoFG7pUjhX3hOWSmlxN8oKOZX+IDZdO76B/mT0
JNRtUO7Gki1cERMdiWWP5mefVLCzD6cKKwy1WLFJY8GHVL9+7NjPonjPiXXMW4tA
EmbxZbKBR5c+2dD6v4LEM8lGFCGjxxGogl0OiIwXxKS4hQ4iaCZHAAfkXwYKdB0M
5o32T7K1pkpM+f4qE9zLamKte7Ogjs/55c7IAqh22LeGOn+ooeLBF9KKOL5dvre4
rUqTXPyGiqTW8f16eMWltvI0EFZXnR3TmlUfx/Nzoa6GUCjcA5ZIZzTT+uxXZWKf
J65FLFUlaOLEkUuOfbTudclsRZJPdvdoP4mJIrh7VD+1LcZTbQhoJeB6hrvNp6Ja
NjkYjPaSGCKdJNf8fu38So7HLgj9EN5LfTzkuD2xLj+QWVYXcatbVGq63k1TkIUU
db/2h5Y3nYLGfszZxKTUP1dIeYNkSLJMQpGw61vEsL5XsuUNprqdFOfikGIu20hY
+q0ryMmTEM8i6YHYyQ120hSP6xZMrbizMlYhE9z2/duEuDjq8GeD0Vuo/31bnVb5
FMC47JVoArsSv58P1eOjWwQ45q+4sCbieo/UovpSahwwx/jkqHCP0dO2ukmRoKGI
rSzyT2CbgAun+z7DsPaSRirqZKC1wlcV2nX2KruEJenOvQ0SEemy9bxPtEQ3/sTT
grdrn086fuY3xgmMMo9VxZjBfVZEM4JYPwDs61h4OGCYmrVeB+3v+/QNGi4sa/ii
PlIlOKTrfburRoz1xcARqsErrpjnu1cq6ghjX8zwasMd7ZpxSiH8q5fSouVGig9a
YZ0KFH6OtXtKRkIEO/gKHO1H0CswQXvxWcdRspOcrUaIfJludOPX5lwaKteneWhf
ifiEh2NWwiJ9Rjz0sfdSe0955raFjfyYK7NfQNm3WjTR55A0QG+KMsbpsiKIEfkE
S11bSE1/t+2GqegIRehhtwVn2N6z7ZSieANdaRmRH27kIRnlP5OT6sBL79+OsZ+i
22OVp6MqqMEI/KbzIWtwhEzEzSC+TsqhshQpw0kQjYqeZhHmPwFH8nF0N+P+0qUb
FBfjxOrEH31wvyTPqUWM8//d9aP8lyu+dxjNfJlxAgunopqeDitHDHIK+nnC44Pa
4Gn58yh0xbLKBfFJiNQa2EM8Gckri6gr5E2n36jQuD/FlKZFtroh1PPQvLJAHLs9
SGblrGQlHLnrHBRqtYYIvkph0Foj6etFXS1io88UwMMmQNMEYB/DEHo4/2jTzcBj
0E1sni3GAYxGjh7yEhDQEEGpmVUTa1TpdmHyC7dC/dabeATC8CDSVxKR2Qh3geon
lPidb2/gjKOA/A+5xIsVPItoL4WC4Y0aQBnzPwHx9/VOl2AivTCKOTjq9dsRh10G
4iaDoCL60WrI/cdJf3EMzCnC5alIuju9CXf8TNNntBq7DmKA5eNHOhmOh58VozjO
1/UhKeuq4i9ZRmVqj1vN//wqYBuFu4neRaLGH7MofaQQap8K2LfrUsGMvkNB4pNj
VZWTjeE4v1QVe9ftEWvVaKErHScH8+9nlxljGlkoL5cWqUR76BQE7TJ0JKKcm+tJ
4CwpL0GJPjG5c7ty3Lq87gzzOrLk8nLbKd2TcUWbpDp3a2zNbMSm2H3BheDLWKGY
4BtKwnzgMvz2fLLRN2oUp683hL2GPOmVW37ET6buoMq3ksu49iQRntG1PwMT3984
+5PNTMRef1myJyp3qrjC6r6s1b2fv31lyIF4wAMD1RlbKuspY1wb/NDVI4RP6Gik
54ESH8qHhCXd9LiRMgHBYCtRX8rKtMeo1USkA7Js2IY83+lEDhz/AM5gOD3uSJ8z
EWTLJvWQFnxQl5512paVgP8UFtoSA8H0NDwYoQJf6EkqW9ueqZph6Qiz7qbrL7CB
Jzea1MJNkMy+Sc32DsDPhj3evXxFPYJHxIpGDMbcrhXHjd8gYrU4jEPo2/1XBsyz
81XLaE8EzbWw2qJtLI1Bcayh5TGtycdMmMCiXJzTmqS8c9IIMD85mMidlQwboYyG
VrQjLjd77IX/rylNNMaLB+18IWJ15LkaJp34oljqB/6nAi0wnTLt07xC0mvoCXR7
jPKJKQf3PyXLbA3mklx3QVXbrFTiJ9IEvfgwjoxehkjF2CGG8uMgQUhgi4zis5jq
PDDcEPl/JoTfpYqWel+BRTCNaSVxcCzlwvBWlq9e1oGO5re+rWMfUzmaFsIOystu
4SzQfmuorCbg1r6J/SLExhqB4H59EAMMayI15jOQQXvyw5TDQXlTbIa50T4KbOUU
WcJpEedPg4eU7h9ssDWBVEZrqx2Y1CJVH5WH6VJ1RQhjmaM39yyuVFm54QPhYhjJ
ZEun9uwpZqF5oWHwZUACnYJyObMIGrTmjg6r1SVaRAwfGFKCiVI9W46pdrwIYpli
zaMG7VE49cdo2QgPxzFOU9TKvYTjv/yrkK48DPpElNHnOkZ6UehYdqXEp9Z5LJCs
Fg0ctkWQI6lIcrTSAeXDzm4y/FW1ElBcwvxBhOkCYNZeLQ7/1FQKrXNuIu3UHrPO
ZkFWwrzJf+IuVtFcFxhougLWcuG14I2pmajfUAUmuOHsdCyH2oXPDPrYOlcHS52c
tiTeHMOq6qpGhnZG6yTLtPCOjrQ4vDGCv6IVuhF8EaTsrLma1LqRcWmzwEB7Vt03
py5tZO0aCQceJ1E511Pd9x0fEXxvn1FmUroa6Ht8QpIn57qSSFgWmso8SjQt0bXX
h4nqOs/K2V0zNc14C/lodUZ+L467U0EDIQRPGfdcwX9SOTjco+qmBLwgiWp0peqo
7A0UT17OKcul0MkrBkgdolxaB9uw0TU1uIKuIiRDKVypKgetFBhvZ22pS8VloKWZ
BtrNKt6xN9YEgwNWZqIMkS8itPrKhD4j3BUoji1HW+3s2BWJxvDr7OLf+8W+HJNf
R6PjbffamZ6JBGtkRiNBlGLC3eA5UcGNpSRmFGU1F7DzPr8LW6RCs55DKsvREim9
e6qNlaekAc2NoPlra9bL56r7Hxc6GWK1hO2ZX0YVLmAzZxqHpkqdQz1c1lNl0zgw
/pD2dCkT6zg7EeEblffmEn7yyG1VZeDKSM4JJuNrcSTDBLh8r1gQsGFi9tRvwqJd
WThU15joAvsayv1g9is3XZPOdbnsB+RDlB4VQmiPHl6mjj2vId0ZTnbMp5QWCNaz
u3ov0FcoY8jd26OI/kLTTRW2nEun5lEW2Cy0xlvkJMIs+2t7PvIwuMi9dsu0lEYD
jMoXXg506qrLJ/U6LgS7EsYdoXDUXnd1e5+F4mZVFsO3mzHywnfMi3m6V4fqMAX6
Go1gob9Lp0+Jj/f156noNxAOlEbzuOSMmhUi11h5zbi8xLoF2/EdM0MpD7tGOLxD
GAZDUahrWzyikaPsYJ6hpOyW6msKFQ07wZR8WmZbyHPwh584rHegg3iUVSLRsQBH
bOBCQ5VyXiNY3c9deOJTcSJL721PpNpCIqM33Ni0W4KINMFh8U/tguDB0T4pwFe+
yS5fR27SP9NrhVlOgHkhyv/1dnp/+ISL4nljqIY5gx67ceM0YnktlSkrRstpangj
gkpkpECV3YC15crhtX6ODgJljxAjOUnJ1BjW43CMqmcyhNauTekfP817KgSPQzEN
MOnXD0GdrqyY/tHBxojtbAwS9TrXGvXaB+ERzuXC3RhDZqGP86McsO9a4lYkI17G
/j34HCtQ5OJiP7aLwG+VcoRDUePsC7aKcxQ1pwGakI4atifBJjECjHoQwU5Xs6j2
9IyxjjCF5xgTv0TYmc2/JRRZ4Y5Eaf44VtqgI32b2vOvQnJBS3N26BmoVOhHIJeN
T+idzoDldPSh+bUnsJLTZmOOyej3+mX0my0rdHblZ8O3ah7JB41t63YkxlJRBjiW
ioShaYu/VZcGztWvkoVsLVqOI1JmB1xrROeH4VZl1izlmZ/oZ6w8GsuJmMXsck96
S/boECnkOItEzQFb7OFUsBITLnW9eFph1XqkbkqRZlUgFZM4AgaSsAtKlg+1si2K
F9nSDUQGs0NLKFofs4psgyT5zjh4CgqYsyFW/u5lSh850Rv0DDq0iMHyEF3QbEWO
nLPVzel0iHkkZi7YwCWfOOhacb1Pmc1mTCy/BKsJC2kjW2AAGuxFP0cXozUhFEig
nYstcj6Rp/bmXSQ7HRGY2rPVxuDUrlJMdZR9rdzDn/Dl5yh8Sv5gyqrposzH4+vY
VJ6c19Cz9QDbw6fEaQ1NNr8BqKws0sae8gSbumpokuY9nDMdLIjBfdaeqZGYL3PP
xDUSOSJYYnD+lfZHcVN1CtH7hzGl/76+gZGD+YIh2n0jZsivM6Ty4JLlflezEXzR
9LtFF4pfwzngbjmP0dYMuD5IjrTO4WvM8nKzNGrmmwQVZUYUyD8zjytkA+St89sD
SOLEkWs+9tTU96qnkfKV8DCaRdXDbQl0Y97W9LfFqtf/B5TbMlZj3QOg9IfLYCnf
fUDkKuUYHdE1ZmyDzARQOWHggtwMXIRiPB6s2Z56If57zoYeUn41zUaZAk6I+mHW
EfDW0/u/gzYh3AkBxWVkZlrul1scFRTEd09Hk7F/nks3JybInTZ6gFvEwkgd3SRZ
mrqBmUFGhzSi8It7OKyHzqK32Yl0cY5izN2ImT+tMjHdpVp1hGY6xM3JLdOFXNF1
2MZOUwd42ruyv4Oz8ORlTOXeszcRyL65yp990XQpYc5zo2/zulPW4owpUqkMZpBV
+NlanXG3C4MuAoYQ3+H9NaBZ8Fvn9aPh2uzYK16LDbzhGiR1WrAUIbeepRs4FG/J
6sOQ50Aj1zwbofI+JPzNNPOP+DMrtb2Ra1lo0Ln8p0Y6tATdMmKzkfLaNO/Uslhw
vNMpexohcekeNmOeXoF9UMqSQoZi810W0LNRV9KKe860YLOQTv0KUkKNeoOy9oWt
/cNwTVge3Dxb1k7LrU+BNznoWgiogwzLixrcoKsj3fj7KbaKPBRyxGe445mD5zwv
VFoEn4Zr0D3NLgjlv/0LyKyBRLqeiC6eRqCPCvm3WRbaemmXwSWJuRvEGW4trJgM
vtKwX93mYf1oDOVocWSwUHDZ+2hxrOPN990BhKvxB3hBsCZXT2PRFHKzRrQxnAnJ
dwN6eWgb8cxUwVDbo2bYCfRAGFufrd/TRPUWZeAPBBGxNZ6U59N8QRDSJog7LOxJ
AZFgXDpGwEp+Y24tFnEgOfnMGP1KR46zODwhoEFQUZ1xjMIJ7uf1EGOqCO18NXdm
XzaxdjbK5E9+nlYF4bnBeRDNpJZq40piJS2BAdnmeOcDIPUEGyunppvKnBAGCAOS
Mu252ZBGVnvPNf2IZGYGY+0xOrZ6EzbVZcFjp1rMRyiArin8MG/w3Ch6EXq9pgMK
Jud6HezpmJ8SDshd7xGSPwgcsa/HrEpQPddg90FK07ptlMIMcyMl5bPW5u1X9zpL
yTLVpahlf7UaNmfz7JC01peQNlfcBAfdEk7Cq3CAOU+DH4f3QHl9Jt+drND/HPXm
PckSl34psCBVt+aBVG5lXu5SxNBUqN+fVS+DdBwEU1/7GrbBoUtph7bCc+pj8vkU
zMicXI9mhbWEbm3dUyjf7mAzhymw/3p8ooBhZKVLRvLQiwfuKo3XQJ0VI3dCFn+c
gtIab8uQLGrQDbnX++57wjElAYjR1v3z8b5YL+5/SJveICexy+mEzCgZQdRRFFjM
RP6R8dRwuehkKptwHUoTk5RQmLfvxQqdN/0XqSkJ/5hn0MzChPlQb8HHdKeH5R3v
s2dDNvQ+xWGAOrSuRfEaeMpw8EgV+Bip2P5qJ9QKev5tUZm3DlZ/WjD4ebzUzlnK
MuEVUyr5Q2gb1GH5Z82REbk0QY1RbP1itbdz3shjmANRpjGmYLNM+9+0LhXrc1WS
5fQ1F4yVIKehs0EVaXnpEzYqUMw9RWxByLCvXYp3TDEJMG92Oc0PpiAOrnJyGXsN
pn2biS56vTBfOMpxzHdARP83D72JJcMZB9Xex+gIO9Uk62p77o0bey89X3zRq9MQ
8ecdd38Zb+RxRTJY1bppf8sc6cpwqddGwt+dj+BN9P9vuzQryi3Vn96Pc/J36Bxo
WGj6La5xljeHuQ2fKIJJ9+VEZX5At4dz3WI5IlMjFCAXg7EZzpffaEOM9FOXNApL
DHPx9AoFFX9VFVaBM/kiJuIxUxXPeovaf9AsiApwoDwRw7Mapxzi9diCL6qnJ3GK
pBnSHwChr2zn3nl6/TnCAVVWAlg5UIj+s7OxoEi1op0ohnsEntPXPdrGLtAxzmxL
jLqTvy7/5s2qwtFZVvOSezYTRZxlbmnV4/4E1Hir8QQ+b1XYDvQNBIDru+0s0Yxs
tU1OuQocSwmTuwUAQ9hmQuPUZz0mAY162/c9flvyVOjfNNw0MenQ+V3ZsXXQGsJ4
+rrC+zfy9/eodYcFn70SnH9gAyekxZwMt/elxmEWCMHN6QPU8g7rnL9i7zcqMDbx
gYsfs50e5BRNuHYdwwZTZ0zw7KtGYbexalU7h9GbjsgHQwxm0bFSVJFuU60xNPPp
r5UfcnSJvyUrCh/3b75PW+VNFMSZ3NuYkpJ9I/fG1P0kPbyOLWiZYBn8RMl+yqAm
zhGfu+oQ3H2AQlxubtFrfduJfqMYfyXynTHXp9gsC2K8qqzVxeqPhRAPqdA0xRft
e5r3yKl/LQJpnhowM74TSfR9aBb4emd7vcABFyiVnxvr12VcFGiSI+C2kcVDAW1s
ayM7ouQGT/bXosWBR05CPcWPhyW0Pzl+hAt13oBTkqRORIPad8vYZ1QYVMxsFL3X
NdsjDj2SMBgEfh+wz+rsWjYKREQVgTFb24HPHaIotXkU6cktMIcg6DRI04x+ys3/
V+gBltvQuNiJsobvNiFFRjVXwSxmod0DCNiidhY+nxHPJmwuRwTpCiK9TKz3I0Pn
msGUMEq0Ewx919KIrdMiuh+PwaubqH10j8fKu/KKqYenpxiditv7Kz6VMZ19gF5A
heKpnVJ4d6iYLwrPlwlJGyt9lg3D6sZ8abRFbsq5ATNbx3z5DTNm00q5iXUR1Tdv
djdGLQdhSUtDDdpEGCoiFwPpmAId0Ht3urEU12CPzCsdmmtokdDilxPrSPvEX4bu
CfyYL22HWkIV0I6rhYigdGiyjJVvQHDVUdLCjdMBUc2h/SdizYI6CNWT6i67dx57
xLOboecFf5y+GDFGk23rEAUxsv1D4a9OFcxIap86gb8Wl4vIVU/3+36Uh7AKoKi1
Fzxtv7P60gD7wqnJ53nTM0204S5WyzHZV4KTn1TL2TJn/u0wlRLrenrRxTGfF3mW
D/ARRp/3saRs6zzwMoAagEaTGcJmcZQ/L4JHEp2PoYRCVwyYhoUiOAsNyUctzjr5
mQZfGJ2Bp47sdRqbXTRmtHHmzWRzr9poHpNqimldv5zlen2VEVL7MgLZOErgL8yW
eZ4A/+Mhm4gGIuX6JjzPb8poT1oO44zFA/bY+DzReZGBRYHmz4sEGX/dOz5w21e1
f6/Hwcyl290V24jqgS1elDAGo44F311Ompp5BHpSHkWsV/FjOspZDrigftMA5Vve
79CjsJtxwc1gT5KCQx1MI9ng4ApW4nR3HcXkDGDYofgT0c7UTVWRL9cPcZtsDPgk
W75e1NNu2yN/vl5Z5OeqJAKCByn1FQmpiqsoWaxR8YDEY7ZqeL7/icWTRTTm8Drm
VfZEV3WP7THzUYyDln1dyJy1XR3MKWa+LLx63SDo4amX6wfgavPEufiIyA73Ja1d
rqoPLbNMGl8sqkJk64Qt9LLtHrIJ0GmgWxVi4u7Sp3APQ47OtgYZ3i46bo2XY+7D
2VSLLY+MXYFB1Am74Wu98m0CTqHbbksy5spSdjCOcetD1zl8FpH5nVjwAb1E7/7r
+3uetEoKF/LPIs2riYtMX4wn4p0ntWiuz52KFSmZaSTwaGa9NJzaenthr4+h11IZ
KG1wt9zVqU0HYMnBTWU6tk6BqeOnh/AcKHV2+Wll++xjGKLUj2/bHUvk8r65Urr4
PKg/iBU08+W8fD4/n6YaaNib1VCfSa+n08VFJEGV3uW+N6BwipecTkSrp7JL1LRP
JtrwxhPCICcNmbv//vcUOZ4MFgpltA5dx9CVYSOcD3nbrYJUZ5FmqFsH+TVFclwN
EQN6sfV32r05Hbvm2wRiRD8pf6+Zbygc2mXkIBSENA4RWDFb7hnCnAO/TDoKBr+6
9JQm8DRhtLvXwCrFRDIXp2usvoAs9rZyrQJR7CAVsDLjQjm3nbr28g/RRl8rR5fi
4q1+CeDrjFE5s20tEfPYQwcJxvq3l6k8DtzK7sAj1ybCNuEEsA42QTJ/ddX58SnG
rPkqssguxHfccGSEUsr/eXvOua81QVS+iaShGr7wV8TnLAcBf/2vj7WmQZtY/jao
74jvwAuSVDap4ZyF2ys66F1i0h2pLq5k6m+/QcBP8IYMoD88Nph4iM6LQLQXG8gk
PbOgJmfRP5bfatnGiH3QO1lhPx/G47mvMk4Vsz6jweRTNaCZXoqCXXbHD/aH8J4f
+CEWOee5Y5TJ5D/gxINRNngz4xyBpvpfaFF4bO+64fXWZAiwiaAKofrxqTgCSRry
1cFWvYi3wVRU7bzvwVx+z3aMFHP+kbE6js3C/HxPtAmtq1FdrLovziuGv1NsCncy
VrhsEYMB3uj2LIQm2KZK1QJbYT6Zzoci1XRkrHX0AT0nz7vrJUQDq5kDgtl8j7VZ
V5WrCwJNDo5AIc7sY3QDuAx/k9aEgMAlVNuy2EjDONisCUy+mnTzKJHIxaia18RI
GLIgkX9+ZLfbLY2/E7LlTDWPCiXzlqOvwhYCnmRhC4up/QWAUDkcBbmoovReSkgn
zil4W7NHz871ku1PxnF4u3NU4EKHHpo5apyAlP3FknVQjjMq+0n8KB7ynPUALjw8
Pibo1ZzXGdWeKLnKEPNJJRO4q7EtL5BOXXiZw5bWXOSB+RrbTFNb//ytm462AXgx
BoFfASGvh6zK3vKSBQ7S88t+g2BAO9E1/25G6EEMzBjofR2PccSkX6glmmIweGi0
R32nIJOxqDak9BESgmb/7yxtPoZMGG2kiP3PgZ9l8mjJwwEf8pvb6ooX0hTXLgIG
eP3qUoqNpyXUYAa9FUSK3RpGGR+kPvgezO51VN+/Jdokf0a9iVclvv3FxyGxeeY4
62qOotXg8Rt52gfOGVeJS3X+je1U94A6XyXGoT3S+trmErEDLkVcCs4XT0mQsM13
OV84uFOFgDKhNATFOBBxVTflmeBLbvVe7Ycdin5ijsOz9C1VnfdwtcISir9VooRj
MeaYQjeuHDNcwIi86K57ImqFdieGWXrW10Wn9o1tIaEaxohCx+tfWE/2RKBjTQvL
54BEouk9M6SaeepS2YeZonkJkG8PpZEvkgiUGiO5BZ1a8v+CWM06WlMWy08aobZ3
7u8bB/CbSMrCOFy0AmSSNiRqWVK9qaOjQKyPk2dQNztjGnX8qDgbj1SiAD1RlpEE
SY5S3mTSJNVjQsIJsMxVtkY1YKzSXF/+2v8OL5MJC6dte8XpAGseku8Zz3J0J8kt
QzEGq3L6gwVD+5zRGD2nTALOMbMcxJJMgGUiLdWJb8mFNwRvBBaEW+e6Ns12uF2e
QSvgS46BxKthX3UyvWXNpuv3ChovadN6m5Fsc9JIA16qBqX/Sv4Lb+Utzx3XKE8V
597slVDGTh9Tnf9KYpAIFOfNU5Fw0rx5e+z8MNXx6ZesGhFykGUJMvw6/wST0lyC
U7NDx9MymCvacLAEPyAyM4BedFE3I3NshEHSzk71cWMasdNFQUqd3jBumLq0LEv0
LgOw9+sNIiFFIRHllmzajp+KFPVEscPEZXBeLkFrTax0ZOBxmm23m+M4W95UHZD1
P9UKiAihGjUGlgZc2QdiX8rOBL/g3LxupwZIa/wLsnuPPlSdRWzr/oaeUv0ZyKF+
VNRa0h7oQjp1tv+4tYW8ySSZVa6JPvdaOVCDg439yvy0sSurCLZMx1Wv307l2t7l
gh/0UttezGoTaUIBVImtkiFjYtaM6RgImbJnZKCbjqO43VHFjc954FZxUDCXRyfu
LDCBGkQo27/OnjmgETDxHMbxdEc4gW8ZF+AWp9FR24imVA0in57sjLb/Te30a976
i4dunnU5mVVq7S7WuDy0D3VUEmgmEipVKGdnfP1XUFCOMua2e8eWKOdnkE0Um/9e
SWS7339Ta9H1GxlwvzgxOGnURcS8qxrbCMobrqHSdGQ+Pzyir7DNkmXCCd1YU/bO
+58nfjqGbyckCcqvKZQwlEPXDF8iKdtYt8k7X8w5AnqtDBvftNOzoNPgFBMW5nle
aeC87kMXnrflDO25Q+iPg646Ev2gjuadsgxfe5rRnU++vgJ31f6Ui9nlxcAWr/S2
oVk/9WRjc4mC/2d29A8yqG/18hdlp68fbY31xVSMiOf8xyUg2lLTHR5mAhaWpx0G
fdyeesatnpBaRRXuFXuM3LTXjbZamjupl2ZkJoTs/RdoT3eNwepeBTj9VwOeYZPn
d/4h4yGTV+FmIXRu5KhZy0g282jsHE4cq49K1dY9COX+6EhINoN8lkDJu5pK2Q63
tN3Mpvsa3wuja23ewjrfOL5uk9TWIXnUkDYCX5aihTyElppx8wkbMBBwtdq0MvLu
+awE95CC3Ebo61Jr9KxvMiWuNcSA/7iyb8XJv1WJGRB/qllaAsQmV/BQKhOsmrng
iQQ8ZBTs/mpuUQg0NqZCL2zgEZhrNxiybRxPNd3pM7EFirdJ75p9D+LZuqW8yi0Q
xRCbJ2/uRxN9a91FFZqlhZ3j35N7WWJsfENjIIjo2DGuEARYXX9+UzcRofoCIZis
g0zsw1dJ5s6AshEyQWOefqET2vW/rnvypvljZM5ds2rgzPR6hhXEe41XrpAKdFxY
SJdTf2bNyC2NnChlQjZMx/VNtx0mLbMgrpvcp9gJbjcPc9v2Dbe60gWJ2LyLoSgo
gVouEhn+OKJTE+kVix9PxAU8XU+U7ZisaZRB7VnfixvQHm7pessbocoK5vtFmHXv
7WN6qXm6TPcevbnGCIQSNdFGzeCdGXEiOuyfoe0bMqMD1CCQTN+/DVSaB4SETkg0
pXCXdlb64hu1+j3M4l0zvqlDFtvf/9gBNiIvqh7rvSYeJObX4D4KULKddiKRktEC
5/gQeP39yPXd5QPN4kIHUO8g6t7gZxd0wTICGMr+OCO73HVyNY5bU7DA9GN8IX+X
NjDiyJkNf5+4UjvaLr2+c71rmPLPPqOd9tiucCwg/03R+BaB4O+LFr9Q+lSyMYNh
IJ5ytK7HIgvG+8PvlQt93dDt+JC/rMhyAeQPCU6j4vL0nKUdanfxQrgz9TwALg+q
Kit499OTpJNuFAXZWGj45Q95HVMKe0MsfMeRtaS4aEARaPy+jU/Diwajdhw/Bj6c
+3hMiOPguI/rR9IsOHWWMt5Rw5Xl3v4DBmDKNvKyAyNO4twZ8XptWRLzBaet5CA5
tC+BB/uas013CUqHxNpWIh86d/EccHnoRaTcXZC9BXHgOMmb5bPAELNqKtEwYNuL
4eX6ZmEPe1DKd4meqnxTwcDrMhd8+gZC9XJQlF4nrXmKjodmbKKG2arbGONKxYK5
XoPAiD2FQLNFGovk9/xVQ0zfwHjY3Q49jCS5Uk+/gj5w5YHdp2z8KHR6sAH4QMNP
L6U8vpCi6gYcxxoZMX+6/boZ08Q7+8sdZPakWIWk1k5WEX+gMt2O89mZhNstHwc8
YsxieP4W1E+UgdK7MVLckqUYz960Q2ob05CiKyoP88GS/KcL17Yr6zdjoiuZRCfb
Tux1mpQX+2+nJGIqkaWfR/2aweJb8xcl2ri01Ong/OTMOzgoC5rvcnvePjuscenf
0NsR2MWPBIyQqKtZD5074sXjFZKngfzQrlkVeDAcvpbGERUNwJ+4jcbi/FREhkW0
UF3P6aUYOFUcgymZ5MEDigU1VmQFiP60Nlm8JbTm6W78CMcBbcpE+sO0gPLM3T/N
zrF5w7ia7fzfaLQPLgt4XTocHZXno6EW7y3dhDQ8eL3UCvrDIGdf1VHml4GWxm3O
ASaiLEiTD39Gnw++09iXhPqlEtdeW+JazwvGT0Y80swynGMCoGeOhHTnVdfPpxP+
SphxDykh5NiJ2itZkc60O7KKyYBLG46i2PopPj6BmTESvHBRRSyBGd4brscDniSh
ht1Nb/5Q4KrDWqRAC34Yg01GKEa9N4XPZ5TBi+yYx9QpRSraE0+fAbyZ/l4GjN+I
1mGBEebSB4Kdj58O49KC+WH7T7hldqzoKMY/3ZxuahJSC5VqHD6+Jd7CVxefg1bk
VE31PHSbUyA4vL7Mv2avB5TpPBFU0L5XUzEMcoyOthqQHdD8zAhwYlS2ob0yuAhu
EHWA63fvGmGdet5Ur3DIrInc5BNe2nO/8zGH+BgGDS8w3kF+SOsnIcEfesqSjql0
HFr690N21EH+yf8B3VN8ytQ4oS6QmJ9QMKBEepcL3YxDSbxobOzkeVpo9228Q6Qq
jn+2ipTonhCYsMMtabj7Syx1IBxwxQhUJF4uBCOQKEJyqUtiXzf8MLQHxcoS4u8Z
isvKYQxra/kirTdm/wvCwicUD3CXXCcdK6+17JZdggJCL+t4XJsypZyYHHareVmf
wcvC282vwAh5dv8jCbFH2c/VX+kWO8GJ9AQjegf+D4brgaB+iDwoa0yh8tH0RakP
mRwOGEMGLaN+SamBiY3LQvoU6z1SBTTUXrYasTcJdureAXRTqeqhnrJrwGlbgUeU
cdiqwm3dZCp9UZ75W1sc1tnL27AUwu4S5IUxm/XoiLEcGPUWXMOvGV4b+Uro0Eqs
kwzBTSh6eKAJ6tiV5qV0qUs9vluu+umpZeKKXtE5w/WLNKh1ld/F7LqMIJWzXTrT
3SjuOVJPkRmfu9LgR5CzrAEIx4ohCQz1Sw7hbSywhCd6LMNG0iosFXFKdgz9HNPY
vjLFvGdp8AxadMseXl/XuYJ+My5CfyHnrRN6iq+G0Aqqa/KjZGn0CYTpd/29F1Bm
cQn1o7AI3qran0RgDPKInDb2gLH/MqG6js0DjjLCyGCKcjiaMuRE0G++VdjPC1DO
IoXmH/lr+dCsFz1uAtFcS5KktMV8UtJpG6c2LqTl3hqZE8/ir1YLEIbs0p0f8zDY
iokJNB1TvCsbtZATNLmB3SO8wsiQSX8Z4vJv3gSS+gZ4UB5K9b/JTvIqOVjwAYdo
AnqE03W7DfgDLhNyrDVk1SmO0XCbHbG5epxc3/R6j7PsHJMVFd41hjSMz+AOhB5k
h6DnbYTPv3l41joeT9KLMh4ckFSXJGVw6LWEVgAF+uliU7GA4ofmDT4XLVaX3YwA
8l/Dr7Ov7+YbstjSnHQse8r2gLhMeZP/cd++S6YbCQk/SyO80U4XDOs0K4rRFom+
QBjfyt3z4vPYrE7gDksQNuSa22TbWPbQJaNvR1YOE2rzaYVW2xT3YBuhnm2Zzv1q
bzuLp5yvQP64vOoB6E23WjUkDOmStGhwt9/8UhXm1FsHY8Tpb/8OAwma0hP+0niu
4ynPe3VL8gCm2i6N+fxSLGKyhlB2O6Zx0UnKGLyLEPLz00dDC/kUkJfvLDieEfC5
Gvbqu2MItmyK6c8dwISCsCxmYVb8Daiw3mbzXUSH2JP3wgsOII1gNdYsq6uKuVjS
nhpFFEJuBSbjz51KPfaaRgvnjxzbYeC39saDYA2JGaXJj/GOWogIcLc3uztm37Fr
jxAn7HUdCB3Ayb97u5S2ZgrvW+zX9Miit3HG5FbKT1dTgK6cwgNPVqiCtFWV4mVv
a5AvYTXVXgbQdgzAEcIQcetySXX+398o9BvYA9Jtft8bY1r7A0yBcBAkNwuA02Er
AzqqfkFTihKgdiVdB4JDaRQnRbWbtnw7nZTh+VZ6YpA/iBvCMUdlXDqNdoKHYn07
aX/FMJrLC/mmiKqmnJ+xP7X3hHKoQPyn6rUxcLHqNu+yGcf44F0AuIzx+2TXW1V8
zhg/3lCOhaIcHwBDoQts00w2BkDT1ez+jVtlyxh9RhKPAkbLFydOCXD8sD3F83X1
7QyPlXguOJmfU9OCZUdcTjNp8n6GuIWzcPjSdyhG4OcTFz7/9NUtbW6VHzlOJIKJ
ObGo+paD5ZwSKKI3W+/qKbppkDely+n/CcEIOCKCiH+de6V4Ehkfw6ijdDSvijrM
6eFJF5plBUQNYCevyVoMVvXfsVlG5VE36ZdBieLECS8c7M2qVBpoifA+WDasId8c
Eu3+62nn5/EFyfDomVLPNTA0I8Ltea3M+5miHcFSc62FVgz9FP9HLViT//nMCBNq
y4CX9OUiHj/FEYOPKD6MGBTgKQaJ8ygoVBFWgNzEJPQQ+KMkiUrgFndnQ29i7P/A
eP3ffo9dzLINxgoTCIOzn5jwQQZ1+Xx4dCQhYMJ4VKLnvdGvhgfkyacREPbIwYP4
Q/37RMn+z2ot54ba8G2fYGR+jVwlz7CPbpcYlaU41ziU9D5CUus4NHvi3uAc9732
+WvwI/RliDr7c7OPwifMzj2SOZ1x3g8wXf6WI0a416vnWJBCgnNtctUyQVlvcQyK
dcrZwcddpo8gLUWmkFJRtN/lBueLTRKNVf3NE3XnCWF/+ISU34OACFEiR3PK/YGB
/tdqLxxYJxVmTXc5NOUR4SHKk7fn/G8S92r7CNNUvAkvgglnDnfcf+EBf/7/8naz
01M74VMzWAN/sbZnVeoxsSW4n+w3K8r432r+BOChCFXgLaRiWQ3AroMAh+2i/zqX
WxwOlQDSFJdoq37koqa/H6f7P6A6qILhTbEPNZi/dMwrqZ0ESOZfxBLN14/X2k28
0cOF+EOvI7odGDkLnV0ZE8mS5VEbsdkP+UBziwXNT42Ev8GdtHrpomeNpCdvlVEw
25tplLbQNWVy/8k22OO1wCg62MW3Pjm+h/4MjGBBPRCowAwKqG2mJAM3RFWZH0EG
Iq9G/AiJEiDMuMHT+HwbiRkE21rEM37e3HoHKPPuaTgsvmc86eRuj/i9ub+LI37H
aNTzcpFf/d8aqnv4gTAeQH+9pcXqIRVco6VLlvWwYXD9By5+8+HIhhQUJtB2CWAz
EArj0gGtRBtrygALZBR8bIo0wyj2X0KUNlLD+OeU6RAYEKwzSOJIOCEQVTHqP6DS
U7QsjIMmZc/qS96m7eNj9jX0IzGIpcb2Kj5h3NmtavYOUMzXsHjx4FOhmc4aFJAU
/x7EvmzyGrafI8ms7wSl64RiyekVyOa421lRKKRZXp3XTPTL3BH26e3t2mM1zIQT
1rdy2uvD4HnrmEHQHfu4OsrWT+quBXbxZ3D2DXzC9UK9HXu9o0uQMU8iAnM84r/r
JFh8dm0NTqfiNapQm+GDUWCaQ2HzqYop5+5B6MsYmIiqoiRBEGStBtE5tewUxwPT
BoHTKvYmX+dEb8QiGdPC+oNe7fb2i8FuEP/WkLKsqeMzfZTRWZ3HaHHg1beMBch6
Z/59Z4dmCcO5oKSNOEIcpmrvYlY/jsQ7yjia+awUh8l2IO9c/w9TUPUConIGLai2
Wfxs4jBC6F81Kt1ffxCzte/8q2v0a5jQ2CuBPrFfL9Wlere2RSuu9pYYtTJrFlDU
muxtcPvFNV+lGS0YVvIKghqYKhVANaG80gY5NI6iI7vAJaG0zH+iOER8FEydKmYo
OlxyhEqv4B8pnMu/W19fFikr/3bGG95kfSIHRa47Lnt0aT3WulASn3E7C4p+JNf0
E4X3A7w/wNHHhEjQnV9w2ydR9NU7SnF9NwJ2u/gygwhx61geUFVaBTsxGUZPVcva
u/HWRUQ9nGSdG9nbmcWNZmMxJELc/QpV5Lmq2ZoS2kqVNqeaiUyTp0sJ1z+mm2K5
7m85pq5mWV1AC5xrXzmwYo5NzvwslcWAT8kOvASEBBBlfxaMCIX7yNp+eBOhb9qk
1NEYC8pFNKcxEERVM2aQTqqmkh0VJL2BXsiIkjUn21Q59wgSg8Qvg0oz4ucdYwAw
y+WEB+V2r1yHmAXYiUUuH/1y7Bb8rOmECMS/oepY8+86q4QAni7xtceYIJXsnMmo
ge20qEelkl+dYru4w1+M43If5nrTg0rXLduSW0+n3RxCA9rE/B4etPAoEZ0fJ3vm
EzKsyDM1xROcA1Z9anL14nj+u9gkFA9mIp9XjMwqCfzNvQ5wKCA8ujF5wnQARqfh
YOgG9j9duyEQ1cENvo4sL5B3RcBlWtDQ78xiDMl0GVBcDWAZxt7kY1Ffjca4DE49
R1owLtdXy4/Gt5yh4cG7YdbW3fF6KN41f1E02yRLQ2GusbPn+hjPeGT8oKKKRzeR
1t6LB+dgJfsirddiOlXw0NQDc8dAZ72ju1dqu5dS0IbCmvI3XAAXRWay984zDvy5
9kA1tmnev5dLBYZ4fH1Iaw5a9x5H0BQDELyI9tdD9/SmfZ+qFQnQiL+m78gADkNm
WaBBnsA6yUfNZALG3Y0mZpN0xAtT4e16e2pIQmsUolFeI5w9L0HQjnI/ATt7J2Xb
E21nfhVH9sCn8lf0CIS/Elev6VUIJcCVyyXH7Ws6nNAWNyFFBEes0v/8WFiEDfZh
VxkXh2yxhA1i/sWZM8uSGHbW2eeFb6EHAY8gMuo89wFZ56RndAzBWaeaUYmh4ART
/4lEuVxiNd0Vz7s6TDy3vgsQyEveZETVeqw0Nnx8y31G3YtqHRqUe5SAf10egamS
UBxym4F/p3GhpL6kIyG2JnoxHbL8DCJnao62b05KUQPiWMq/02tg8aEwy3ULJN+L
p1JFmj0mOKkWqlwgrZw3NgZjw4VjfsKmMtuXZUvWVU/0RCZ40YTk4aJWnz3dlgNP
5kMl6qkmdTNXte84P1HTZgRuhRHCTDYphL9oULry07DnLhlNjcuyUDLRMQODMcpX
o2oDGEMLVbcI6zo0gTXHCn7pfGNbXdtezIh3gzpF+shayzicXBUY1kOxBuZvIiRL
3C3x4IVRacfnkFVcTzcqfNTiDaqG2L1HdIu0uvAZ9TUq2wEqIrMniZWbXUdUAi1T
LsSvTHkDTBwJXfubZ3RCZPYdhCJY7WgleKU+xDVR6+3P4xa8k+CfAo+6T6X/Dazj
TWZEbnoz+DhFrJuPixUPCN0Mdn8ktDedh22egUCfUGAVx/xO84AbwPqSHJ2uVJWT
jBAX/vrg9VGqjeI0Tet46F/pIUQXEhITdAmPsSzk+N5yXDY5jSxTq2Im2rzFSyx0
lk0F4dK2RixZ9qjGzfIbD8Xh0CJfJHuRLmEWGBbGWrT+nDft5EQgvEUqdPPWEGHQ
I1SqXBKdg9P3Oklbo6ExQWdNiKDLSzdgaUyASHVds9J3Kr2UBwf0ZVsO7sAxBV4U
QzJ5UBw8k/tQY4PNw/lAW7OAN668bI1qceZwJr4Awv/DanBvua1L3BLTBKLoFV4d
/S8Qy/Dh2e8TNpcG+hBny2xwKHPLQWykDQgOlM7PiTuLimgJGVgtngUW9k2bt50D
5V/ewzxfGR9eq1QzPaMTJz19RSgp+3FHdzwta+2zuhlocJQZws7QuIZwTvZsVeEc
wQbN05f/ZoYRseWS+C7GnlsBGT5WQzg6+nzYckez+Bt9HlUtevEa3QiAIIWkKtzj
IMUSmut2RO/2fbFfMDwhfrh5itd7UpLToBq1wMKEhv2S6LEtikdfj8nhx3OEj/96
/mBwxcwAMdaaNbsaP+bMzkVz6O4SCkbkTTUUfc3hKwmNouWG0tJ6QbBvN5nzrznz
2LfYGdtPn6/LufhbhVa+oKML9V1iFzEpnF6kigaqpHO4ochJVWILgE2rwa0fbEO5
jumCZ3vPmaGMvHIA/wDw9KoTVkxM3hfcLWjylLg5TBcXlJ0V1jyOt4R34HTaWl0A
tHYoWcYElDmfRiGbXP3dlnu14H0TjrSUcAzVbaR3vyPjzKJb6qG6qu5kSsw22yFU
gUVJOvloINi4qHN6BW36j17w29/WZqRcCmebrnA4C16iTFORIGVxNb7JeGaprc2U
wXuwVmroIBjwUUIFLZXe1FwrnlPO6NeuqBBXnwOljTvjRhiHR3un8HLHxLh/t3rN
kWDwo3mwRwHG6AWVDD92eKOVN3WxaCB2RK8jcYcXNXWhzPJNL+Qq2+ciiGuQVDJn
DNbqIForJvrlLJ9rxtAzP/CbugnqpFLhS/bOXJN9Jml4x62vrG+ocPOt/4ZFgjTi
graNAgbtX7RRgzXVC6atWiliWdl8RiF1tk6wKAo6WjLm9JB2sYzIDXA0M6kincLO
uQlMoNRE5FNNJVMEIRF8FR13FKiW4Wep+4ZCDAj1fRNf6ohAVBiPuzPHnucAdD0R
g28f/wwb6nq7yb+LXJt2wqQ+2invX+aOgCfcDOLrPNo9+s1LeixI1Re2sCCOxqQS
JHQuLHZtCgiB+IDtaGbxo+tCBS/SaPOhTqjzJ+CRYvd/fXd24rJk+mp59Icg1LEW
DqNZX+kiCdY+iduhSRKpH2JJHf7MsWhsqtiugT0KFAGe/wRHPodB1kGKwR2fDH2I
uOojmy9lfctRDwRXXEZIQYCAHwVraPomEIF2ruGiomyhNzyWN0bQn3RKdXIH6K9m
gcuRtRaKShBzflrx41sLLr3xqRPk9qnEmIIk821vN8fMrsSZ/EMIkX3s8b18IajM
TftAfAhR7RTPyqdriWB/foyhYLswBLHIKvidLO3Wjva9uKjO86gczNG9RgEenGJ6
toG2Ldm+5sKo3C0xNCDOadhTYbbVQTGSKcNRU66+5NUzMFiIJQ/TCgVZ10i6DDRl
BFQiLuMWZ3TwC29+vvEW1rtZEqUdrubf4eczfwAGnpmqHaN8EZwvInXXqlgD8uaQ
rkvvVu7l9k2MGbVDvaDMoa2+dI3sQ29Vo7EuyTC5g20EnKWmEcD2wzjdxhOkELyM
X2jl141PHrEpgqLZAFg8navCQr7UASwFfauF3p7KsX0DLsfMOc86KRfOm5Gf8FfL
PhCDgUvswrufiQoHqeUFUM4o0Tj3wG2s+VbOXpsL4E4znnd61cdbgv42ivr5KKih
tVhbfQ9692p2p47UYGStfETcB2pXbISp7KvYhPJNlq2HRh2ssQrSjgriXIl8khGX
arDWWrUj7X43hqGfhb3HQq1CMQKrSbfmeea6aKzdTq8PGOon97SBEXKbhLnULOyl
g24g5b+oLZFuNO3jouOzellnaYjxNyncMofpYLUBaHktGH0LXNFJNYbLi5ih93FP
boOhEUlgtiBL/l/OpG8NZHLgHEjY8aW+O3hrarSv5iI8EqM2iJPEC1aRKSxJ3vGt
/KgXApcC8SK6YDlpYVapJ+zrN7bm6COkj6z08d5euq2brZYNvDyvJ+DsFafwTvMa
262Smml1PkUw4B1lVV91LDHKCrrjkhwxquRd64G9q7m/HMGe4k7M0/fD7fIt49D+
8C9oFW8efOvit9RjIFS99ILrW9gysyHpcxTjy9ObjaF1QxH+cKAwqCh8AnXEgXqf
HtEpNfzJE4anmY82YetTYFyKitsFzclSTkCwEtlmhzjKDRWH+veMauaninOgqSSk
cNnkMAtmFNxjV4KrLD1WHuCmxNUOlEMVK2K/hm06Jw7FR12VPitGZ68mDbBV5E9K
inBXmxb2Gohhe97LUKMOMFAP7Hso9fURQsKZtzWv49IIZPlnYx77JIPHAG20x+2y
36nybXDQICfmdEwVxp1akaCd4h376MZo29lSwHH9XnFNTqRIpb40iwO3aVEuoJKs
lZqhMMI9+gInRUqKsWob9ETqGmWsPnKFEIYqbY/Q1RfGgpalu9tcJXDgjngRaJ2t
QGZVqbHFoBsIfGZr6BKPaf8drtd+VRkzxpcGYR40ZLfUbX+pvHyOsF9aGjvT2Mwk
DqbCkHySLuOO8jD8BYdzZuYIPGnO/nk+iwhbcuGiUgP0kBLs2thYt4l7s+bJOMsx
35mVGV04XHcc7ZNYZT+pfq+KuqN9f/NFGtQi9Jk6wAQWZfpAUjWEWRXoRfFnTm5e
DkUpKXjSLmR0hKCYskFv3itTgsjmXOk6Cjj5AfX8JVON4Q9qtJvKX722OEgUCXdc
pO0XjnXXobFMIs9yVLkCi+gIp0MCVjYH2+UhB6IvJu9IaidAV5bI96scAsKYaaAr
TmpD3gThuvqj9ngeD/D46W7lG9rRIIrKRJXEUleACoWk3/ML/cRaygKk9V1AlQeH
JVK2gwWeLWDNwmivmbK9+fgq4Ll03ucBmEOOa3WEP/GgbOcDQcP5ytQ9AMovDu2k
nyCN+uKKm7L2CEbm02ECPlBC1z7i12+DGE/VhE6jX4uYMPNpd4mPuiscEsZ1+haV
JIesdqL2MlYTsmH8j83ktsbtkd5pxTZQeislZt7jBJh42Tr6NR/6EFa+q3NRnO5D
cT9tdn96LYbpVSJzKMGbbj8HU1dGo7iL6EM5iP0yxT/9enIGc7x6LBSza3muYPCb
2Iq/bjfB96C6smW1Ajr2D7JCKMh12s4+95YWBkHdTTjObTsitm7duDAl5MQ8EYP3
UZKgdo7zCCTaCVt18bxGqI9JLrjL2ZSI2Rjyqan52WaP6r+aJNWHHb36KoVe52f2
x5COAXYnHG2EfRBvyByXvzfEj37Ijj9LW58gkGjsdTBXBD/tnbA7tXH6uDuuJx0J
b3ukAycpIMSKr/iIKOmDObxHVle6E0Kyn6/C3kvhPBzKGXLwV1bxRrblv9BymCYt
56WrrhGXNuV/YxiBXjMsR6KAw9d5yGh/F4iqA+Sq54udGwo8WLNROChbOeyangbq
G4soIqz+igSyZ9P1ur35yILFUJQcDz9JhcM/jtKUCwJlwJTjGitVAZRH0EJA4w7w
vk13BFdErP8nfOg46TsSPgAfu/q7iGnhDG4b1fqOzxcKf4YxEKmyK5ZTE1IveWE5
2iekg86Wa4bgOCOVIIZMbja3ZgEs1IQfgvcExYMmqOb24zznqJivGhBsrVWxaMdX
BLuLjv3lJ/6hCDBi02tZjy8gq0Lu4D9Ho07gx7iB6kphjapMVwRR0Jf/6b52hlt6
1rh1t3me2QiJozrphfvsn+sAfwopIfrbuor00qEnM9NiZDjojSjNApZuwHxgaqMJ
S6JJ0QijvvpfQVCuWW52UCa9SwUGWIWFKGt67sIhKBvbmP2D+IfHPEIcCy0cMxDP
Iz/5M0S4wAHGX1PMHfuk1dLPMo8Xwdds8m9wHfy97Gs+XYZzRgOTaJzmLLU5Fgcy
ya1S1lo2a5fOohhEGy2ZoNBdkKeg/XZ1PNoSnvDuqk08r0hTtXKMB+mgbJJM82me
S99+vyrD45UTCI8vd1ynUhdCrBO8XKV5GMEZTsd7HMvyW5fpqjIYNvFqLsN+o4yW
BRRwEcvfjeTveb9EDzdzwPddWNQ6LhydpxL8iCNTmkzW/S31hcg4PZ2dRHWBR4FP
NQqaKh9hCRGfIIwLjTBqjACTi8TwVGLmH9SiuRWNlwQdtlp/QhTyTh6MZX8ZMWd/
cbMBHPi0eIWSNiADxWsp+zo+4IUETNSzYBsuOaDUNqp0DWszGd3gggNQsAhGe8FB
ugbOMK7PSKutrfnGpCsjdSNKV32Cuk/9sTUMuZqbESS0OeV7lVAjNkexY4DJFB6o
CzwnhsNQYuvUk3ypXXxbAMt6IPTAQ1CWk9l6J7S/As8RCiLatgRfUJD8ZFFmiGGt
UpCVgCdr4h847PQbbpXSbh7dbB4xffuVBmIhzctk/s4Yrr/+gvJRj1jHM7mctaY3
gqMneNruDXppFXDVtZQX3Hl+1aEelvms3AzjGtVGMlnVWzAFAh5spUupM4h4eOLq
6ONms2yOTNmJIpRdvARqGh0DFt4AdJgqRF6u2os8MxOLgOMuAM9+CpE+pnor/sIV
2AyccO2gFweh62qcE0pzyJe+FNfvfE6RW3wrPz8O0UYE4zgcD1tZP1LagKBeytQn
rgABIIbzbShSwr6yVRe+veS5+JbzBaVboCVPO0CCYpCoPvO1uqMOEAiZednO/zsp
uVVkA6vpilAwTo9RZsobfg/CN0QLWw0otZMOoFgiuwo3qenHKTgAqCjTp8ZLlGtD
ZKRRcQAGViUEG4zjzUYf8OLTde2vMl4d053halTXmk/iKTTxm6MggP0OkaiKGVXq
O8fhOc+ljKxvGEx09hKUR+f3Zf9ITxe9E5O89U8emBqF0GQyw/M7F59EzFUWntiQ
3SD4Crq5KqmxdDp9KikgK08DRloLoMqxQUmnteP5FvEMWbVaqttX3lUtbkxUZx7O
qM7lUdD3NLWFcOBSOYRrWO1ZxR3EZMVcDm3ftMfFiRnLWlRl42ydNrYG3GwpkKdS
ReEv4nEbC3qt80ZGLHgF/SvCK8stE+lcBc0gUMR373NepLMnEVCxgfAbAjljJ22R
unFm5ifVFtBDbb8eXaZ7M65cwAj8oLW44djW1otdQf6EV1g7jcd//zs/nasTHXC+
fAtagD1N6jH2fQ/s+tyStG+GQNdMMPdQandyOmdiNgiFrLHTRnY2YBrx+AD71YXb
doeF5FWpsacPQdO838uQVgKqKdaYIdXiZdZ8bcpOMLSWDsZyulPhzgWiJzR4dIV6
0WieynkSFj45Pv8CIgI+eOPy+KFSDBidr+QYxy7ywhR4yI5x9GZRHQdr4t48PRas
5yQ4GWYSlL+HMsOy7r03sWR/GNFmmR/dbVU885l6eDHaJiflE9UKzMDSq8eHuy6u
6qPUHwRBc9ECIVDA+ciJTA+X6IVkJiKVyhEGqR0n4F4vEt5ByMHygOWqOc8/r5vk
3tOxBHxISIU7qY8IekXXvqdOqD4TlSEAArGQIE8j6mxy7C8fv5SJej8+C/86j5o7
uNfhQVla6mBT/4d+cRfbC7GqHiKWhPW+oDxJqVRDI6+4wHybovc8YbvbZPWfXD5H
NiwbRItAYglw5kpYIA2R0cRH6DL598s7cEuu2umHNNEbCSv8OEz65qYtepQD/iRV
3dr3+udH8fgfNxGFSuMMl3iPJpPx68lXLb2FahANejkwTLKvfF+/6xQhN+XSONP+
F5frlNeizSjsHCybljVyrpi2Pwvgbii7OmdyG/ydq+PYspjUw7h5uNy1k86RRNXf
wAAs9X2eICXIpDS6QDCiCweiGe5o7Kzxh9PYCjajSP8ocRONnkt2bBHDqqJlQI1P
ZmiUnzDXEoHyZNqC31Jnx1Eq4+FLg0OHGLfz45MQ6CiLQQY2dVEqoXjoSi4LLd2j
N9EmnLsasu1yb04Dj3yuyW438VC5J9ZlIx2gfp/XFOnkVw/SV5n4gh6HhIfEJGVQ
qEv+ERvyLbFXr4PPPdS4YCJCgSNW90lmptNnJDvkTuvnYBpZRW7O4snXwrpf7oVC
Z2npOEQNRlHDqXVY/8YEsfDWAIYc5TOrOEyuqAkYaA7AWB6nJZO5eF/Jl7yhaV4e
sZb97ErAxvKSahG1K20GTguEnQgZLhSoL42bmmSLL/817WRZE8eNZVSmqHbQaWsU
+e5kvl3rO36E/UTxkFsn5TugOz7pqmTAwLkDbG9ry0/V2AsVcgXx9X8cFiUsNpqi
bWVDiWCJKnUTI3VZtiyky3tdQTFRNMa2Qr8FCOaZjWXDXIyOIn9g/x6ErT299DZD
vRFgqSnAUUj//WWizGSGLyTPXfgDyVvrbvANzjPrsolaJ3zPHHQFzl2Y1OwALSQU
29pY1MzyvPAALvogXfwjolTrMMiKGHR/8AMCSxxQIQpjZwGP1O7o8IctFL8H25G5
B/osh/sJ9qOYF4ihnqifUuVXcgF/MZx4n8UWRZgaFWna67lQ/T6uCVajF3Vrmelw
R52QU5R339J9a6G6LEkOXTo1ehrXSC4W9rL74lZ97x7+UF9e0GTdMNzo/MiphibI
FJVaNeNtMk7gnlVCdAWSZbuq2+1eq3iSt+eEptt/vHohodmWbpuIhxGMQtuAvC0c
5gBKGR1rw0NqAt6y/3yHlOsHkEyrPYev9dNLN/uQWzL2SQ2FT7VybxRZcELudg6w
W3CIrlZotfasIytnpUlcKkXX3a7nF0O3nHYe8ZnkJ0lx5u+ryNhYhKLQNouejG0Y
1wxwpThuJ8zxiUD5oGcqEuuUVGAjQfwdqP0zbjn9MgTZ5Cuq/L3fp0mNwn7jNYkv
m0PVJbwZZToeYLqDOxug/m8qhm2zQEWLXZpEkiF9DNWcXFSUNyGB6kKdAdMaNG4J
Ps3EvZ0u+0/41Sk02vDTBtgjLqGwznocYQ0vlng1/MQ+jOJd4/rmyfWWKvhKqCIj
rT7JXa3oWY3HkuwBI0T4P+VJHZL8HhtltbioOZjbRonhn1nRRjKrF8/SpaWr7bss
4ihLach6WLVWKXsrR72cziMGVeCBgXBF5p+zb+BvdnP04+CAOxMjhlqnMNXnKSR7
JG8HpuXmIMpnxde6A/T8tijwOD+dW22QOcoWQs90dzG13IiJf55Juym0EeELla1R
ZXzDavtrLUBgGA6LJCYFR2ufK4bmimJ8fstq3MpZfE8eo/N2Gzl9VEhwrIcB7cte
LlT8R2bo9NTNfL1p5VVPZj4HvIyonGeDTBu5WXlQRS0QYGQvihnWeSgES+nHP8Ue
wcwbJkiH5G+1k7oFz7rxtofgE6az/LpbzKp78fVHVeP8yKvHbRPozNwmg9xEfx5T
MpUDl0Oqo1AO17YEiLXnvE3MkVbTBjI4nul6tJKgXGQUXlUzLnQpYLl2/chPX1i/
58EQxX3OvvYRdZuzLIFV8lx1tMBGjEmaa/BYvF/6fdaZ8imh5k7Eg+W6eMEW+96E
UuefB1jkgDOoZ3+XaJYkA4vysdBttrpqgo4Qs+m/Pezy08VLBHmtcIIPh1FmZ0d7
q1QowVMEGeAJcEP2W2psy6kCL6SVW6POEFBzqfMwIOoC+T4/x+3jDfCc54rSJ9VS
NQ7G9l6o22lkp8E+ZHObAEt9cyWMSTj7PUFTyvbB9HGY4kiw3eaevAtN5fT3OTPF
4jcl0pHeBiJm55fpdF5xudzRPvB1ryGzJpygpWJ/rYe3lL3kC64QICLWFsavaq+4
i6RVbn4T6+6Wn+i6f5Pxgg7YrMescKWzgFqiLnVkNTGzIo+4Ff9sKhHnN2OxEKpc
ScvBM+1QhyL+LJD06nN3vwma8KRnnfZ+lOLVu3DMeUV92roUJs0EJ35nMgELXtxW
qM+TZCUtRZDCmr/M/QadtxHnW2orjKR1RpoCl91vwkLvzLfcCnfdPbP+ncO7g50Q
Ohy+tpvm0OuPiJdS9YecoN6p6vl81CdQTsNq9WXmcV49T5sHLoW71YXGZefzZy9e
/n+wc0e7Pn10Ov2bNLCiUNdWjcskpl0iDrU1Wp78jtzqYnJsXtxhtE0EQGfCEz4K
+obf6eD+jrLJZ7OrFMkBrXissELztb9f6QRIbr20XYwWfonu5f+1UU0z3VZueWKM
VbVhmchO2j09PHpMbaHps6o7VkKU733ffxxoJPKWPfeV+X3CJLl3NAVA6TDyfDOD
zQn62tG8tkBCL4Az4D4c0hvp1KDx2q5wW1oWfQyUPMgshgIH/dV7mAPFUt9mbr5w
YFm0VTpotl61zl2gAdORQLYS9ysSHaV38In/bBXkj7JDjjLVzknDSoSx2G8X8Ouc
5rLKKMEn3XTqahLt6mcaMYLWBI5TW+OmLbnHKxoUlkH7dDzUQXTKYBs8bMtDKFrt
1sCsGDEUSHy9WgNi78yiYHUGbmHvjJFMx5eeS6EBJ9dWXeRT68DBXlWuJYHk3TSH
eUnjzqo6PL+OCUh6AXxayV22ZxsXs6laLkckoeewroPPJjcGOMGfLbrTr+pkg7lT
eu421mSmo0wftAqLTcqyiiCn6mlzsCIJfeP5TgcbxFHn3zXaQQgS8aFts//oorW2
MBdT4JQXDJkcVKFpZNzTU7k2qISTQRisB7FirzysWKq0uP1t8h2KtSjkOhTLftet
V965tWYsz39tQ+CHoSq6CzdK51Xmi3u9mFmB2pXmf5LXCcnkUDJ96JP56vKlAfzB
ZrWE9c8KpCjNxYOT4pQZAafC7vyqpBKwb9dGJJKwW2Lk/sRLG1FrVmX/jMKhgXo0
flOpVK0maVwnf1rOcpctJ5jECcALZRZwVR68PX91Dvy3B7iYls7ZgdAdIgUbV6yb
g3y8tiBMopj84dzwGNxUk2AChHX80HY/VE3G6KT/x6TMoHvzgtYAPW6k1y82gx9R
ivzTxUZpmQRfgG0uQWQoRymajVFir5h5TDGv8yyiQTQRXW7X+Xs2b8hvJY7sK8Xf
5dd/lVyOnHCqGevkQscrxrf4Id4NC0A0ME5U2iOSuNwAl+RWsotmMWsSQxDkHrR+
79AqxXRV27LF95kspotQvrZiqYOt9S1ajDDyONB/qH5bbyJs1Yq1SdzaFSj3DMVn
UPorFJqNyvDaEGexd1TGjsOg7l1RYOpztPOaX8TBfpOeAaZ2ar5n+7wItCbdfOi6
Duge3EzNYooCUYTc0ltoHeYNebzz0p45GoeYtH27qScdMFok5fIPCZUazf1Ts0E0
hXHE1PXyf9QjAw3ly8p6tCXuAK7v/2zvclyapYq652HQ9y8lhX416b6l0hIcpq+S
NllsUShcpCbKVgdr+zTxTUwGitJ0cyhctWy+25i1+KG0Nv+nDhkdwjsDm0l8cwWz
vtdELBhAtmiurVt+llO3cHP38kglai8iWBpXxYJtdb9J7bkuhxX/r8b0vvk9G7AS
aeCKU1Apehda6heYagBU7PTl/UqNLjZniAoNIoQjEqquwc7HnZMtXcRpAToxQvR3
llNZH6oSF4Y5LjPLfA/IaUN2HTqY5pM1rJeEfjPemaZ6SR4jbEuvoi25x1EGhqtl
cvUIzUbZCO8I1vDEqDkmMOM8RvqfDd/c22iTiyU9WhVAxtBbkm1QguOOMUfOC7Wd
BhGcpU2XfPi1258Xv4B+yLvd4twYp6xxJxmGr5rfHRjaSYzN63PTbgbnRE/gcGdS
VIyZZvQtHJ5G6Diykj3i3jhNJLqYYFQ1q9BogXqX8MdiHwmmslRc4dRK0AUc4K9x
o4btBn9BAFrDqnVuzNtDfFgBNOHQnIUV/N8JwaCv14lfkWIrNmw4ebUegNtuIJ/H
0hUy5LO5yAbC+X9bG2qCRZZRG7vomZ8Poa3hgZO30Cafv/MkJyFI4nKssgwYHRvk
DZAzfVwW6BKRS830sTVeim2NLPB5h5tEJKQ06n0B0iFLTXY5HyDYcrsd0010GCqD
1X4MxfC/MVEPstkUAyTNjjmHRhYO3WVTE3ZG5xKF9l5m/odzRc2C8L2GD+pzztd5
FgHHD+Azcew4wRLr1ydscH3+diAsksd/R00TJEqbR425/sNOs0QvO9pkq5QiF85/
zox4hCGn8t2frftZbRXL1M+dHC/qP9GlV51H2mEh20gg/0V1oPCUUeF78+/6Olse
uQMZsPaASydgp92Is1e8wjTLKOGat8sJFGaJZ2GbWy64U5FthkE5B243CZ9CDdJg
a9kIn7uy0Ki09U96dmISU6xqcCjmggNHUmYtlgNGGYuUFPg8iXEbFD9vbOn5eJlJ
9vJRFO8Q7DeNc4cwfbkWaCzPyYzHS8Y8kq++bsVUTNnFsN74vuLrvbRswGTE1UII
U6G7fPxw2a27cw8AQBs/XG3yvx04QhEc+iy+7ychwsb6sqJepeI9wlUsp2ZperUS
mdpi6zbiBAxFG+KKEEzoa84vlb2yp6y6I5g/8hs/dClG0qpATMZJ7m+0PUEnqigA
gyAzMa3/yic2ZJBGdwHcxpw6vnDqSBYVVBqErN8YntoxgBXdxJ83dRmS7ij/qP9J
rj+9e1q7cygAz8sQxG05Aqgtm063SorlDbHEMjgCUyqcAnahrxF7MM+f2DDweBGk
xwhskR1bUlESbdO6NvAXqTtvzFFmONCkBqFj7/EWw+UkwDJQrWfpGFzFJ4GiQHhs
XDHNXG+V+4Kr4RCywyNdS4qPz5yc/rGwy6nksxN0Me2bVJapnJa5KHTQ9tqS32LF
CslVd8DZV89Sn/0jGVRv3pg6pf9g+9AYreH+L8/86dx9xgCbFcNtRCy+TZZNJA65
LZ592ezho35uFr0JzAs5HCFcVaEG4XhtXTldTmG4hJFgkO9MYilDN1KAVOFXsQz+
5Igr6y+zNtHwi3LTofHhwGCOZl+NQEK75i5D5JwZVsDQGA3ls/HuhZ/H5V/coIQN
3Z+7CDGpUoyEK4I7LIBr/VvJxhStsLu9Yg0E9ZHw9mLbJiHQb/ppIxNVnXHHuEq1
X+H5uGzDmWCiVzplIDAN1I8GXXzCQtzSTXKig9de86hUV8rMEtY+zpIQ9ZI0Olw6
W4mfepIaQnym2bD1lr2skGXBQ9WfkWDPWPHQ3Hav1aidTgUBi6CZp0w/JHaNFVLh
e4ehsOYdB0Jm587XIzs8Xp1z2Agcn1VFg0CgwRTb3vmrh75kZ6OZoC+4JPoqq93q
1tIcejcHs8xWF3f7eJQlo8JE9D8/OFC6zEVz+eMAHkq6Zv4iJJvCe9F4Znxo//Fl
fKmRxunT3jw/FEEWtOJnzPmv9G1tkF7P/xt2mtx8nIjB5wG0/So5UgUWymsXl3mg
1q5JQmSPUcC58rmHwcA5K2aVs8CWEWngE1UreMcZaP2RBj05tzKqmwZkBtDuVxbC
Dl9UyMGXEuj6vHOiFtJgZowLEOQyCM1QJFD8FEBxCPfq3vjxGR4+nRbyqvhjF2x2
DInfAIGz5m6+DFdlCNs0tfFy1/dLdUMEkhdyZaXg2+kWL3Jo58S4Ipcuc0uO/f5p
HmLPZKQNzgesrqScvxIjdsODcyn+iwzKrZb2vni64/rRovShLkI/ta1e0TZj35dO
91t06+FustrFJzJ5ljnYDaBIrR+gH99K/E+cTYP4I5lcT7YrSp0gpXBHjIeqNMuW
Q2zHCW6lj6AzChvGdiijsekg2pdz5/EWvnGBKIAP80sHhkFYwxXnwwA/26PJ9vzu
yBYX0k+Oj3JpAozQufueAbBMCQ5A9Eqmrirg+LialBAQUoy8PUs2Bo5F1DfvaMKh
kEG9UPncWgHj9DAeG8kKOm0QPXg8gdLJQzdJ5W9oy2SUsYZ405TiPbgsE0oztVTG
QzqYlj9nKeTMY0c3BcKcTVSOtQrZH7ApFKbtsk12HfBMw8BCbJDth4tGpgH968jB
U6pqbzvozJQ9SsV88PQ3cSvm3BP3k69kQBpd3T7q1dXKZA/Ln9f0BVWNxcXu4IZO
DEyYVodaKo2PclJSEpekOWtG3EVJKFVVHK9tF+HZpJnhp1WbdHK7h5fqzNbJMt0V
lp2ESTjBi4vC1MaKI/hDVhDLYqMYXUXsVuAuRru2EYOapWeXyf7oH4dCKy0t4rdT
zZH3Wu7vBNdJAbz1OHi/sVH7hcm64bTTaOh4uviLiR7YGFXy3ybbPPECRpQ5i0og
nr+OLQLo5fIDKhkGvHusEv3qRn6u12G3mUCVSn5BoxtvzvfUHhMN6S/NwDw53SnB
VdoCk4ug5XOXGgZu0lNzdCqb3y9Z7Df7mj1ZkG0ZE1xT6OzZMvT4x3OVhW3b3Bi2
O11XYnyGeQTaTAygfgiq0m/kXCJ2vX0bCv7NpUHs7cRnDw+hypGhnH1dGe6EMVGC
hpxJSaWVXfygW4a9NaZ4byG/Jj8MBPUYIOiyFXmP1moRYSLEHkJOdz+DFWGDVBVo
CjyqRjXycFDMFuHScov6RZhy9p9G1aAJLTyJpgOiGMPH8VZ39hYzOl0CUrCcW8qe
k+bByqZBzAjmk7Qk5REzTaZ55AOo4YIDibGlVFRblH1uNgt+ZlNjzgKeeQUkc8GQ
i6BdVNz8ek8THrcliIG/TXmcOi1JQnlULU4+M+mviudjzVrdZQ6XfrueCl1zApZ3
tXJxFP1UK+Dr0Z04oVKvPmiYit4WDguylfQHT7zYNsKQ225K0Zmu6PSHZyLwveYN
8AGwaFo50l4Sy/0ZcbCpISg4jO+yJsDAnByEcbNwBcFLSB2oK4X/3f2jIesegHeI
Tjq6NMcGuigaNcEoCKhAZc3XyGZ58n8slQXRNckdbKbjbbxXux2ahLYUjiaVcz57
jU4bioxAU/WiZ8bQRhtwPVC7I8/cByRofe2hiBF+VsdDenvG2HUIhjnvJKlMhUuy
IwdtGqTFosOgHiIxl1trsB9IfXYNcJTkKqT9dqPGsZ3S/ez0p3nX56KyNYNMcqJQ
mw9fkmmpy6ai50MiZqcFu6AKAuP9t2G9zUHrZ4IFK16YYBWZAyQ4yRm4nyZY7aNk
MLjZToCb1ufyaLStho9tQXPKXO5ETiXEP9Kfsmtw1vKAVVVoJWwYNAT/WPTLbx7g
K5fKQS5hcLNP+wn70bqjnYRu8C1rQg3IrYIS75p3MBRtUjbkt+UlTdD2RRagtkaa
mXUyTezPuKmZOwRSIjP2vqdL/8NwXPYdlIjEDDdpc2yoodtENFcjCiJB1G39uhKo
l4tUWfJioylootKEdYum0d3lgbLq0mkHAbOC19PHik3t9UmshpwXChkVH2jH21EE
EHFRM6aXIAeekzQSwktkFZULYoUs2YDOwG60/jogS9iNQ27e14YPGjs34mzNRYQ0
AMI+7D0K/UvPeu8AJ2IyORftPVrW8pPz3NbU+68BD/ekKhBr+w5UBzdVgsNghiE3
tD2bFOlo4mPNVdRWM3S4ssQ2RhjXvNDUNdTZzG0iqtSiIBGEW0cPi0rb4RFFK+mE
KV6IrWKKjavYTrV+jKYSq15U2wDZXry/aTNKegHneYUMy/Re1gu+39gdFMckYiQ2
u0KJAxeHh6XrmOEiCrtSE+o0vaBMGzRkPdGTLYmVVwkx9Fn8Sg8ffDaHCzFfLf35
/LxAG78WNXsuWooOH/bvEYGRb2BcBC5lkY7GQrHt+kKkE23woSpqjqYVehQBuCxr
x2DCSi3F4Qz/ZhxybYHb6f9w1k7sv+cPI9LLIBHtuLuqWDu+thcuROIcYN4ATM0J
r5CjRUV08kww8y6KlpQti0gWZ9wfscvgAwKsacHLStkfzhmqOtU7zLnrwJeSb9pi
DUamchj0ThNgN9fRBzXccuCg2VBrmb9XizesqmxWphjTwbSHEsNK9WUtiB1SmHS3
jVgzBg1QPwJbiH6jlMdsWOu78e1RnFYIkryM41zoNjvNX4eyiIL67jtGv7JiH93U
XaR4AqN/8b/91KCOkZ2ZKLnctRGQ8G/iFnzqu+HRbm0MxMkk2ZvRRxW9BnrkyWcC
Fag1DK8nVkRXwCp3L5SSFVpZRIVKgLvpD4CP6YCyVKSVIGEI5u7lyD64KQvZEz9t
GOLHkwntw5iRqu30okFieS9jU8oRgV+W4QPKaMbOXhNYyy3oZwBM1jy2IYuxV6Sj
SPSZISpXNlp65EI6udPVQbAQRRLcQbGj6slnKlomkqZ0CjBV8K/0yV2XHfLsbCxD
kEtHMBdBjshMb5YNVDqDrH+FImudteRYrdwRtaHqJueKXhnELjEvuIBpXimHXMAR
hOMrCeR5FjhbTfM3oOMu4XMv9PsgR7zDIF0BjeszeU8O1gc+zIdmsTYNLH+W7/yX
YrFzB9KiiB48LUcffHnY8/hhCbyPqdyHb/lI6J3Mag1qndFbMpMeqttnTgSDQQZl
jneuIp/KuSPtKZwALzcWUBUsCF87uimW4zaCcLruVBkuYaYNQ/1U8KxhRFY0s9WG
OdD1HMlgmWJgscOYJFBrn0E+hKwTc1QM2Q83mgRET764cpdx+cnjeTGY8UJ0480e
iRpn7M60+/xfkFjwjiQ5d9wpjmI+MXdciE4sXqMSLbLjP5HDmleM5ANi7i0oky7K
wLHz7TUNhhFnr1Fzgf01TwRBtnA+kfy7mzUF7vsfvi+8d54TB5K9j4TH4FKH9d32
kqFguuWAJ7l+1R9qf2jnx7WnNAxVDbVXNCP62I9nG2KfKs647862JBDp636bDLNu
aBM4RtbHb7yJJy2V+/vXzxToSkFcdsHRvk55Bos7eW3oK/Ya0Vib2rOEZga7NQsF
z6f4ws2eTTZknqvK7XByKrKKH3Ia2dFKAdSvp7lDz/Mn/yaKZCW1TXDv141rCEaU
I+gxAA5Ob0Z2bvMx17E43Ye/5oeJBb9r8CTNZF2yW1wpx+Jj42DXKDO59SFtq029
BGKPJAghP/IBxW1S1Pd5qDeAmwHXn9DFMmEMBzOvciX+PJqWkSHVzjQQak4BCg72
uboq7rBzoBNVKJDiDz0GR3gUD55JYXAUih3HBHtsUMWfH5MZl1KLz+RJBwFGunzV
604cUDXV5T+GS0hanrHWqnlb/vUphrkBZ32/YbzBbT0jV9hILARD9GcSccSeLfxV
cyIKJ1s1uzGY226TKNjR1g542+4xl9RWxB4w7zlYIxv+hqT2eRrYj4BzHLbQKqvP
FcsYGezWGFrUpD4HWtKZyNdlZLzo9UZ/hmIa5GH0ACAlRQ90x0bLgUMldijjyh7R
hchnDhhVUGP4nneAYBbzwLW5xQuBKuXgay/Zn3tdmdDzjO+JIGw8cvX5ZolessUm
tpXddCuvWHJl2TLDfcL8CfNGmKmNs0+7ks1A97JU5yUadq6CVr6I+6u7XmF+vMJ+
W5S2XpHgL1M1TWKyE0A7Q6G3yOetPjsnFSEJ89n5v7ppqkvg+t6OOJtTC24bGgOi
JGHmswsUIAB9LoQIEa0uN0YkKZdjUd43MgVpRp8nhr+1XT4QPtQoEBeVwH/h6Ndx
/h/HDPw3EWeMUEhKSaty+5vbNcKxkKb1+enXkjkDYcUGuabKKpbkoTAAGFYAtzX3
W5Dc3kT5qPRZrnVgGfiq/okz5k5buEkwHbyWLpmabSBTJ2cOEtTV9AXGFZVIwU6V
cgPM3XsCRpb9eRWtUt8OYblmJV6MwfjIp6wO9Q9OVdyAsmjtbkUjUQeR/r05AnZ4
T+L5Hh/a/oI+hc+FMTUjZcVXLLAy231UoqJlHNSFJtDveykY36cciwyH8qn2O/h6
B1tRiXVLdq0j2idAQut3YbAGVIYMPAgfebl1WAI/p9W15Ek1nKk+JDT+cKsJPmpy
uQsp0G/+X8EWjHzh1IBFWEfTRbHBgQK2s4SKU6Va455Tid5xmte1mMruL+SV2H62
Bwd0CURQrrdUQNn0vqH1ChUa/tRn7cplnJtVarOeEpjvG0U6YaIA7Ua0AGLlexHR
XsRHhyqIZBQM4MnK7GUPfo9ujJiR6VbYn/G/9zPOcMGcC49v7SRgCCkIu415xtFr
jV55C8rbwlehCaq+MVx1KDN+Z0GTEIZNDG2iCO+BHnjaI7h8I93CSfiZ1TQsoo6t
zKjZTjtWuaLNJhIEMScIcEDNsv/uo6dXU9QEin0Ee8kKH4Ww7i0lCMgZJU/eR9Bb
jdfZ4HEuyflY34djfuj6Vj8fGt8Yh30CN3+B2tkgAGOcnGNBUI/8oJtivMRJ7swU
WcyHybxX94OyxeCEP6P5LbEDrzov/lJ5UbNCuGCYhOXjMALv8dZvK2VkmqnwYqhV
mlva3q4DpGzCON0PU6iYhshx0ycXf5lk0wamzuUnuiKkZ7RRoxPA3/FK7DEMmCkW
VqxS9/mlkgS+Mmsb6rQIUeQiE81pEqe7Q4Kg+JlOaDMlzi9WdTXmX1aj9vavfIVb
EiaEA+64wsDeLJdh2jIqWUpHfINg7e+ep/hA3ORzS8mTfmevkCYU2EEnNguJ/qC7
/0tBW1C4ERugQPLsrw2P1uR5K+PFQsMQFjdkjOYZrNWL9qhZl0C3s28BvAljQ328
u+JrHRkpCfvEYpj+AYCfk+N8rsg3K770DzJ/UN02wlTJHF+C4fagRv6w3l8C8W0Z
6CfVCZ/I0NW+BB8rddHCwHtSPZm3lwJ8N/32h0CxWnX3YNDnRwT+Twnd3t5y8xma
IXKiihS1nY+C+COzOblkOpM3bsaYT94XU/YPk+iw/f0bBTxJ4CUB9A2sIJ9KO5Oz
rye4cw/eSH1b0/LXOgjeW/60EPDNtjCzunD0Lb+o7GaBm0Gyt+1FuQ38w9Pik4dg
XHaekSvrDoPdCJAt8qx9qPQ1W1UJsH4976PEDuBSqoawjOE7T2CAzHuaGNeULmLT
XndjcLWuWfQOxWl96m5MFm001xk0kfEpjvLVsqcmv3EWEhq5VTQf9ZKBrZs4YBJX
8MGwR3URdC+68jPh1ICHzMcbCb0HNS1TmxzNJW1+GuSDiIihLLAFmSqSiOpgTkYQ
UWkHj+2nXoAuKvOLNI+/uwYqB5laqWjV8Ti3WZnPOTAH8CElfxTiNOhWhgRXO+Fe
fcrkSFVcQVRHwTpcNPJ48zGWwliaCpjXKLZYywh9Y2SQ8hW8fl37MoH3F5GlFJG2
pX3wiZXgO1NGBPB4/ovyctx2CccPq9dHjh7b1faxNsI2WXEpJMcz8j0qvVxE8xir
8895IJ1e7rTnpqi/iyCkami/19CpXvQGjqeuNKbXVY2SlOfKn7VsBkmytufj61hZ
WeWyPw4koRGWV+/+GRFX31KB806Z7blw5RQGjirX1pDC4x5IwOAq/9j9AztN4iD3
3TPxHWC3tP0NZq0Q7Q1cKhCnKGK3y5+4UiNrAmaaF2VCdTvVjSt7ZIBO2G5yUc3y
g0AlCJJYP4De8aitv+6DAz3QGszPY9RYftxjPsUC4JFVo7UTXo5G+TXWkAY4PORC
DQKimTBnow0iV8nfWAyyR3ffQ55kG0a5djknoLX7F3IhDnRUk7DVXPcxobiH1fm7
iKDhuTk5GeudgKAG09+uxJbzTAW4nZyhx2w/66KmhPduL4zs4NnhgxqYLShTiITl
xqIv0xy05VmtPZMoKkFNbMbUvRjCD4FrG7KK55Xzt8aLaqRiFY7U5Vl5IPJKcRUy
Xzl+cW+TtCGEIeM0P03MGIiKEZBqaQv+Cy3SinCD2fruUqWGxSFaMsxHWsOD5EMy
mEC+bBsMqJIVaBIhPWVVgbxrRtS8fF1UJBZFHRBw4RwMfoNbk7MnC8qndfX0bMkk
xkzJrdlZkRMlDP/czf6B5fqeXa2whHgFeizcKk38o+PPXkjEyuXWuB0DFcV8uVk2
fs8+31VYYEHqmBDoa6ePGdDAht2HjW12cy93OsMTWZ5duPY9RuxM7HWqmuMyQAm2
yN5KAN8xG2MNpGXwXP6DjdTu0WimRP6y5hF1SY1UT4QFYsyLjOySgg4nBo2/Hqac
0j9RMblsNO0ed7L3q/EhEfiwmcSnhsRpS8fm7rqpTZVh3ii20oFRYw/GrI/m6UEw
Mrcm5K0oHJYbATmZ5+v8s1ic/AI3pGV1prYF5vzzxvKJH3SF369o0M4s4f2uIlLi
p0r2jeRxzrj4A9n/O7YWVYgEpyTbkiqaz4eLBVsyA7vukoKpqfHxPbGLfWETn+e0
w4yPLR84rDc41VvP8WQfv0rIToMTFH/mTy9dW9JegBXF7wXtcJgNNpyRl58YFRaz
UC1OtdYEYDzc0XKaSAAE4uj+y0TWZj/0+IVnZ5j1Nmv85sC1lHXnL/0oBrNesfT9
AEwKumQHn+NUjON8ystDuvyZYYN1H0h0oZ4ibw+xjOM12RYZTOSgYGig9p9VYgsj
h3DOQ8oqcFYSgf2GwozVLYhl6bOzdsVeCS+m7h2mKdb9RJNByiUdCbi+ekz/mb+Y
pucw6oouCxyf63udRfjktnbCRCPfD5Twzo7K/zVWiTYwLH85oR+APchJ2bpZaUpV
1fAjkNWxzV5KMKNICtAO/gPKOuauWZLlvOP8ZHyIrQbjSAh4WVAjmF+aMcNWTRMx
QRFtaXKz57BGuiWPGxlijTsS72AL2vNUdEwLX9E+UMv0CB/oIZc4XvbED6wXiHmb
9kXGBsa9Qka9gnzkY93dPogA97EAOdNNhWNbafuXt0Oq/BzvZXmdfup37H4xvNCD
z3zVppC5kP1Bmcx5yU7DcxDslCJKWp5w6QBHw2y6Xn9Y+8IRr3f7LWaDjvTHyIst
PThArlaxyL/JO+KggFi4ZaibZ1CE+WvbHE1ixtysVworyQN40XbwYxAQCG0h7JNB
tnwSeVC+LEHQ3x77R8IxxQrhHCx3zHLE3Xqkj/PxNDte0+01aA5yADyWtEZp/+Ds
xJWRjgT/HPgJHrT/QVm42vz+IkqzPD2iJ/gYRxw+kj/D/QsYlbpDe9tv/SEJKKs4
46ZhHYlKTheQ5EDIpX5Krk5BIjsrC1vEwDkxQeY+6eh1QJ9gSPpSZ96Jd7KBgOgQ
rVPZTDCpmmzSNdyNfxXwBoj6Dq3wBNvbwFkH4xkjhFfmg6iphtceVydpyUGh9H+X
QNgQmw3JTLEjVBCWhJHYz/WZyZXJuTZkZMu1EbDlNBC/ngHpMdMQmYBNtfVGevW7
KS4W3ggBE1vsuNPh4HWfHeoWv9qRqD4vWTBYP94V/iUHfIH5lA1Wurdhwxy2sVRz
4oziqTabcmmSvLqczRg4nJ5DqNGy6zcyq3+vPRqZ70F5E+CsSSx0x6B5o71TewRQ
eh6ZF28FxB1IpWxKIQGw56Nu571tQGi5+QyxtqnJe1vpPA+ivPAPFrzx+TcgNsL5
lpIoRYWxrXgfgi6x6HNZeUeGAzr0pHoIL24hGq6Ywe024ZTWZR9PjWOH0AZ1pjUA
ml0A2VWKoPcqtaGHwz2EFBLEzBzu8bH9RQIVJotYoOTpBCw3RozmJBGVix+m5AHw
FVKEsc01bPO4hei8Fh5Vs5qF6CZ9G6j6xM+gWQw8sxmCpySdndEhFr6TM+b5IX3R
qjTO8cOisMLWVXQCHkf4O+rd7X2brPlwIn8/3cjLgE0yqjwuuaROhBAzPMm9EoKJ
TcDVo6uNm5/muO0dmvDEKgIbH7aDEO8DcfmG1iQ5DbbsszypvxNQIPC19V3FlewL
9q8j9ix61HhRtTE+9NNMvCJJhlEyiIujYrl9Pnnw+PDgqQZ0T6CZ8QG65sJeeFlT
OBAu/DKGByOzUAf/wQONn1J1xLkBO42rjtUEjaKd6uFBRTp+MDRBmstyP36kQkTB
4QwhYU+Ruytfu9ti0XzIUPHWKS7IcQL05JATBVOoxiKkzZ/FSz3o5Xle5EHPi4xz
dCzgnJD2Z82N+fXiThU5ur5WlZnSR6FDs55WK2aaKA6Yi/koZp8xWTR3GQIMzBkA
k4j5wQxnDfAW7tf91FzZ6En01NShhRf+DVZBiy8aQoeZs9duyUTcdlwFX1bsRlBX
r5vL2WATKzEeGuP7WyE0KtFD2+WmELmp8OyD3eEyeRIcW+kCqDpehX+DU5iUAXMi
VGZ8UQT6VJGjIMyaDYovCaCg+iDMAg4NQTE0bCCY3KfjxhHFle2+zbbauqZtAEsA
S+zlWFqa/5rAh3fV1tJCuwFyWZMHbckczOvznz9/UXkI9DSQw6d7DfoeOfvwAhUf
XX5sJNGVC6KFTyEvnXPBDARMLa3Otd0RlMGeMVKxPSct4nQifL/2dQXZrIGSO4zm
8KDE7C+gX78YfeJJ8DAkIx665Wld9lxLrvK6biMWbwewporbzqocjLJxn9hcgoBX
a83CvBxUH5aAnoR7PPul8xUH+YXtOI7DEjqN1kflRVknMjoxQMf73JFw92XNAGm3
VIb2avXOgNWocsk63zHVQTE6GutFcAqsrvlIqbr1oSY/zNLF/eoxuGxKu1ksUg32
qdkPdlOn/cOr1qBAVwWKcO8jQx36L+obPjPNEAO+k09tr0SkulnXJguRW6+ejfV6
ov4JaVrW8IBS+9OUz7xK00vzmYuOWmkTHsgT9JJlJPQA5aQ9XlK/G2wOialjGC64
9QPNLjHNDplHGRuhGGZSCzQ2lPPQBgOCeKaf/wRkuL2oPUPrsaB54twWHSiB7MTN
2jOMe0YEWHntTavcTGHaJ6lPF247O2/oNoZXYFpJa9IAESxJiANy1WOwmgFIuzQo
i0lRU0uXfrtcC+1+D3ekqH9/bRPvG6wQB8v9NWIMFPn05vrsqA23w+6wc7vhhFKq
bZza+aNvazMJaIuSIonhHRSj28qogAnBGgaJ2KD56SXBHKz3I2pK/KdDT2b4dkHJ
xWM/zGsl39RPHTf82ZobT8+sErE3uJSJhTmXOCFd7Rv5yrUiSjY0D29YSmABOvxx
OHxZ88PcwndFU7inVy/t7UsRDHqhKjCbuhw2EJ5oaTwBup3mfSL5k8ZkwWDCyDf6
9BhCaXwZmO1O1KLxzzXDq59hJaxvKvHUxIJavI7FQTgVA6UqW3N0ToVvrQzsfZSF
ri/bFotcOBVJVBaqj6rcKPM0pXsSENYVO4bsDVhggin5/5PjQYqxQnvqFOePZnlq
RP+EGWMAKq06o3o3pguiRYL/ztn7+clDwg5QK/9hsLQG0YDztfJGJ8igZzasbVFm
ZHDVrdZo5Xx3N/nb4DjGG8GRXj6BuJ6ErJjKJ+a4aDNjtsh55z7sHanGkKvMUGbX
r38fqqO5MIEihi7p1M63GndWSp5DLRgsQpggpHrNM3ucahDHYJJGeKizM0zWh71l
6R/W3tAOojAHxiSO2j8DBqDg/WnjgA/zmwU5yPKMc8uKzuvN7PVb/Nmp+mKCadxf
qw9BGtKKQOc9RvyS6ZThEIm6xXvyUJS6KblUZSQ6WEPyZkflk1NvgSvZqGpNQZSf
PzsnJfiRHWPGa1V1AF2TeCnunSGwIYHONHUnPRgSYK+a34ZJmUzbv/77SMYiFfGf
qfs7P+B80dwOzO2BpyhiOZdE10JziFHDpkp8zT2bIlth8cOOQ3oerKQEUPMbTwJO
XeYQscfLbZcI78kuYd2HdqSwpUk/iDY4xWAQP9bMILTLMBGm7zquHNPSns/m+gpl
Py4Q3bCVkA9FnfFE3rjYlxgP2wc3VMR5fwYjxLLeJ7xrhs7eIkqQtP8ULg2LOawL
ySVtNBLjO7xNeXiaXHlPmN6CrxVRCQbVe3dSodE5JB+8+oZnKiEizwSfXbhSyCOw
oMzdGYYK8TShd1KvbkoGA0HIp3qolBpB3G17an1ar1Lo+d/ANT/BYS1VQ+3VrtTz
CJraJsOF0cqL6J7TadpJs7JQ06n4jl+upkKWONb2papKQy0ge3CFVKiBsMRWEGuS
im3o+2hCFCDbLozMVDjJu0yvIlh3c4s27R5H/CcklZz/VPNMGUHChA9b4eivw5kE
/NHTw1VYU3hmgKQeNGy50mRET4eh1LcCXJY++jobJXZK+I3tvwqjcReERbwIm0ja
Vt+dMBGkXxLPQheUyW3KjGMgVDoxZvLh47/b7nDXZfdtZf8g//TZ/z/QEBZI87ji
eVPOyof7BB9rX82qH/2YmSkwCEAeeCM6/eslm+ZdXIdagTvfSciPuJyWZ4syXzJP
79gbthE3DlWgZvs3J5t0cjme6BF+8ZgoPfrXaXNmT9GcF1O4QF1DvVux5rCwcztg
Lm5Lt37XfBwqqit0Gvm3ghKK6GGiV2bl/+UvDnFLPZGvADimu8M7PtJNSzIjJKJ0
fldbvrS9em2Ifyv+BpcnJg3iPdeiFORf9x7K5S/FpSRHA32bok++a8KUFSltN4DG
8OZj98AnFbSaqjwFEzG6KfVeAlxRZbUiDYmVguZrYxsLE215kRaqplLnZP4ZdqDr
jGDjDKy70TdnNnJry9MaVIQXIWCBJjMuwOT+IQ7E1e1hiZ2xjN++JLOqpufQ6Lqe
zjx4IjeNK0wrUBv0m+61x5a+ZULGFjeFMi4NzFHMG5MDdw5w34dkr9nqmGrIj6be
Po6xtmqv14+Pw84vXsnUvy6KxfM/UqNcoBM07jQWNAea9LToo/ZiiDWbCI7MOe3C
LsCLvmeUFd3jZz5RqeYcJS8/nQw8dAOxvoC9m7dg9DpzxZsUfn9N5HnBn1lpLYdO
YJzzny2Niz39essq+jRcz888CXSCx708FuNdkFpbcoFY1ZlQiqMh04AVl64X+eUu
MZzPh5sa0r6meM4NivpBzNAyYzRY93Xw6Rvqa3p9b2efz3o4WocbgWr4CbyLgjOp
G+5xj5oelE9hmNbHcb+MbzYrknSrij9t0zPEWV/Z58o+0iQv9JopluhK9NjdHyl8
2IBeEDhqcE2UThgZ+78do/JJeEkrkdPY1nTj7bmc8Cja1NLsp9xU0kiiW+XPTP8X
O4fjkZvFDqjbnJ3JZJdiWTYzjD3j5wurmoDh5cWMNBEGs0HfUBN4aj0ghJ2Fb4N6
tn1L6oVhBnuq7H9ipNaaiu0Wys7sitxRLSw31I4M/ZMeu1ig8W4qPm92n+nCLX9E
bklhCZN0foBhXrAdXksiFqZvVCvFJt2XcZBkO6QUuUNDBK0upPR+KJeWD8VWt2vT
LU7F7iM45sKAgC5mj6PFozRjOOf9M/FvL43y1laYDa7+iVvXx8hwW4NwQY+F8o9w
TDH4HLBUjAiWP+sLyxPi1x4Q2xkqSNk7hIuFC5G7vBEp85K1O1f95YckS/z2mY+Q
azS3NT3DGU0MQ0/3bb/4sTgL8Y4JCC4O2cl9H3yfAJASEADKFPRUjBCxGreFd+Uu
HWFSVcYVw0EXaVZrYI7OQYZnzN3ZUXnL3pVeweM7AzkYZC4FXxfQ/Kt8swwKOFfp
uWKdnXVF44gvdNjsiXqoiGRg2ak82lqRdB0TG1jnWu0qS+fkL9hW3B0+3zHfIZJ7
tqbdIRql+XHUxq+iDHUIekWwhRWJTKB7x7eVwZHixaENV2Jq7jxLqDUyzUV0eDEO
UjNH/YeSoC6gjW+00sgJho5C+gioWDhXlZw3fX5L5sVCW0U8ZjM98+POSDnLqFLD
9LoAICzWFiVgEbj5vCjoGlR8mhinyKx4IwNH2/L/083XH/EgRL1QA1KyEnwCPPNA
nqTPScPaihBB1SAYCEczQRuO3z/5T8aRxjHDSPS2PWGLHD5BiSCV6jl96YvazsXY
FvLPoLYTJhwL61r4skWcIeColGvlPktFdchAJ21/feiTwqBqzzfq66ENB/8AIVbE
UOJl0t7crTCbm1jNh4DScDVE58hTce33qf+14md6klEMhwk2GU7Te75VlXx7buDc
P1tZ1PhU6JoW5y10tGOE4oBa+X9zdmEUkKmtueUsrKDomZsQP8dTyNj4xwAMQRaM
8tu30t3xGKq9JqefiWA8NK2tz8+vOvqFGIn16zrsxA6nHWOVKAClC6uLfEipxZwT
DyMjHy3YIyMGpH91lQp7WTSNgMpcwMfVyfHiUNPLPBNhRPF/Lg7sP6d+71pRbtE4
Zeh4UvCQ3u52ulVLvI14UnCsy2ufaYZbSnLA6MIsFr9UHVVEUTLd0IgS3/CrJtLu
ShBQ+inzFYTqWnuE1sq5+N1oLeOVmsSIfUUGsNMdxR1Vx+rmUfWn2jvNWktEchN8
52q11rx8Fy9v7T7yQngX12LlHKBH2yUpR7ks851xPiEEtQ3MjubjCwqPzUQXbhi8
Fmd6U3iwmiq/0Z9skw/A9PeujWlKOq5sNS1smvVTdyQbClwak47vNLyd9n5xJQnp
siGp9gY0xO5NSNGsHotzzCt+ZLGQqYr1OhgsAb0hskV4S2K8V6wwapyhr/zh/V2g
gLxu8QSa3+u6ixqkzx8J0scBjHRV0Do6ZQ9jY+TMES6lHvq1nAty3l9Zu6PozxLH
o+rKk4MIRVhN6C6OxhRHe2tT0F5w/r1tCFRlDXa/mqIcZslezc5XaNhgdqjyA/ob
t8VmrV363iq3ETUS+7GNG7Sp/Y1TEdQfckYQygZj7Nb8pHDgLEPj7U1VZ7x3u4Zh
0SP9mglL6AnPsq2I0bff9TcWZZdponE9J+z0LuzjVWpGZhAikiUmApplW7P06Yx+
KByw33ZEKbQ517eSpR6/fHP0AU4b6Hm/lKoLYD4sYd6YxxMszQyUVae1+CaficsI
32iT+x0dcVph+iFQS4huW9VqgbD9dT33sKrpORQVdJI9Wl71CGnTwIX16Xc4F+u/
HKv9AJRMnjpJ4SjsJuBJ/fM2ZEJsriBCjACOAVLRMDTmwIWtuuWVDB5Iq7VZCjJi
mU+BS+yXERn5A83w5y5si1P9tWqhrHBrNHS9DmJmGFXmMqVegyI9Rsev+t9Gjplc
OSzFDpoU70yPYC91Pt9/2/p6m8zzfG/pTbKXsxJYbH4sM6ey/YcQgDOiLgDaFzIm
JQrAO4VMqzo4EDmnrD8/H9ro57QmA+YFO9CNkscwKM8KgAVOK9YSFhjV0ZAYiYuw
NxQJKvxNZWofzzbH0zdmoUsRv/6qlM8TUb8WH3l9stHU6hRG6H2OOfLdPvFlFwmi
qPplqQ5AezaISNZnzrOECAJEqY2iYAbwt5KRM8aL0H1zuLnP1TAXXoyNE3jE+hoo
TdgxYl5GqbImoQYSfR6j7N7aBQpEjpBZ6HgjTRrma0nso/oy4Qs5KMuDI/gUA4Z3
KuExijtJXBDIljixccbafuqBWjlAHuM6qtQUW3JL24+i9taxk3w0VWSo2ZXOfVoB
SqTPUW/iHy54c/tXvpaZpiz/I5s25Mpr6PMIfBHCqlcKXlpRUOKiw5Xjml5rhMeh
XmDVyRns8qAaAF9xpdgXr8eHmoAr+pD4bUUc4fFrwlaDuMhzo6rJa0WVifaBQjZg
HR6y1GvZfc9HiK4gRib081Sx8C1wE1DL4wgZcF31BoVlg2XzUbVEJnCaeqCG6CPe
Qr9jmtac44dztY3+NLTUr8jgy8l7oQOpCPi/hwwUbZohkii38QyZc66QNLgRZq22
RM5d3rBddqIJzPPm4sXR8HE5e5aqLkebZn0HhegrEDsDtuUU5RRggAcDCSbO48DM
lh2bLMHqioIWP799+Gg7mYergl4GsJDzxU1Z6t+TCfSvUYPBOvy9/n9w+G0aQ1k3
Pa0Ov3qk208aXGx7tJSO1ev+3hN3V6M1EUM5jmTSQFnamA50HiSpe8Y1SCP9P1zu
RraDAWNc/FA4wKLpaUrEMmx3IzdlB/66Cvfib72bg7AERfTuUusk5fHMTE0bFJ15
8CFC3kH3l1jHNKLH6rcLJOyvWiS7OKqavQc98h9heB2ATxBN19CBwaikzcAZ1Vwy
jIjuavEJra4Pjy+Nd4YEF501OtVjDz9AaqmRbxGoovsRHcA87CcRrJSlM4lUICws
fuf3VSpLUyG3gXgxaoJfYDb58E0jAdTtR/vPyhGY5Fxtd1VHqFUWhfDeeXyyVlqQ
m4+yJisD1L/j9BSjcxrXSMY7KcY3S4IcVtM60OBsA2k3gEcmJS96TVmoBgfdoRg4
cff6ojvn+911nvNEoGgbFl09VXJ5wkv+/L6ex/iqYgz8hMdJ9PAJYHyWxWEyc44x
6AeIg6SH9WrtqSyMiOd9dIyrko4ak0tnzns57nMuVXW0JquHAq6EyRgbtRhDS5YD
YySyVIIOrHPLE1X7q9w0p/+s+vHovZYZhcN7QoYxg21zMecGr8tt6U2bgnHLjEWa
PcgaPsG6Qj0whql0cTZlh0+CDsqDO2N+K5b8kOlgIOUB8KQpjh4zIIn2Fb9gpNpR
TZNZISH/bC5XzC+kZU9FZsBdh2x1B017b9c+TFo0TmDpO/bbHARBr3K/CTnEDYI7
+loTlTGvz6DWHnB507Wu3De4q59XHGkJJR2FdBupNRoqFx0EfLnVb+8Hionp6Cj+
4nVXnvj3YMclRVtSzYS1aw30Y3SkP9OihoZ1so8C65zTjKTfC4DnHKIpzZXseecZ
O28wFwBo09b6uKB1G2egRlmHfcd/Dhl65LmjfZ3N0xV5t8i3r/C12b8oxW1P+i0T
5M9dDT9Zs8HrQjZaELLG/1QM6TETmvyITqu+qPBpS9rX3GEQHYnXRlOEe4KRDVEh
AY9Yk8wi9gV0Q2yKW8AGXY5c/DKYq+qshEl4wbMjsdGJcmPBhH3EvF96t5W8YnhO
EkSoSlLJZUhRCnmAIB2Zb955eT14/8XnW3p8attwMlJv+T4Obw+xnSESjON3xoah
erY4QhWDAVeY1Z2myVX30Auz533Rt+Se6Sv5ITAniXVItT6j5jJ9QS3kkOmU9Q35
bEyW0YEcsyao42H+MNFdBdgfNtClVRW9vdEGaSZ0hebTmgkrDo04bEi9EfYKgesa
sYo1j+GW7nbgXs16fOz3oXa+3Ev5Adhr8/kYXz/IjiU4gyNGnruvB4BGELID3eHN
DPMx7CiVlap+HtZoyI8iPO6DSGTdN1ZVb2ckR+x908QLyN4COlmpozldO6AWGRrZ
fQ3/WHlqgNQh71fSpgv31GZe7AJ3qPafPAnvOrUpAxdWuwVnMf4iTqa27mmFh5pb
hrhtnzMPmWalQ5SQsoQDM2EGFbqldkQaNDHqHpXoV/QRMjRQ8QkAnRJvbMi4RwSb
b6Gw0e24bTC1sXbrKFd/chormalMI4qvThkfcq1vrzcykLpeTiKuCGbcq7SA/afB
1Bh3o5IXezYzHzOJEfrU32p04y7c1sVbkMrrfBuTXzQZwbcCLFEndWhXXJWSjwO+
GPDLwYIW6Ge2oz95+/1RQ8iQMj1nnWfXW6JQ8fPG2wPdWl8J6Bbry4LY+GJUW2G3
ojIBOdVwnfqxbVeBMgC8++vDPA4Ggo6qlE8KkIjuJbLAjnyeSsQXsz7TkCAaL6Cz
/umzXYrHhFd3qEbZKu888h/GKOEi6h9vcnfvsZt0TRo6yV2TefnXC6XTUeAaBs2O
oaHWMO83jW8H6d0m9qU0neqLDIIkUX9IBroJonXwmTxr/PU73rFr5XTaUJxj5fkT
Rp5QNzX4An6VEppU43Kxh7JCVi1kd/ZbkXTyQ8cPipVBxXeGUfc5oK7quSyiHx5V
7jG9zWEBmkJeK7fnNRbojJbPS4G5EiLlfgVtUqZu1vw3h5VIEEps2UrFd4pmYBGV
ZmZOO8uH5gIo1cHjSqC1B6uZthFJg+nBxMg0lcOfq2e62bO2q6/0J6CbVdHUdQfA
Q32l/AStoIekDigpP7pHmlWtPcWKVhFHQZA9iDzKgRpQwtooAiJLL8ev3uuBIz0Z
TWPVAUFPuK0XW85/w2Kl6mR69xx9jsG/XMbr+ZFBH5qbNk0QSJcRRHya6dQfudO9
+kI0bCiTf9CXEya6Ugb/VanEoC3NE5Vq4upw4r9ZCnXfLWZ21eWnopT5VLv8TUIn
RYwiVGmFc5ViRU0jtJRe/4vCyaKfjLlVIdPCxLCcdM3oftfyJygPRc4wiPBA7dIp
4LQhv8ubtWgNoBi0oo1tz1ycCAa4fjAZYe4CzT/kaJWMFIF+O99eCFttlCvHkYPd
Cmj4CuSXg7XqbFrJpVEPX3/hKdZII3F24s1sdOngumlnx3KatRuAAh/WQPOC7mgS
ZE4jXnraF+heq0SgzPPMYTeribRnrUy/RbTvgOQAscYOGEg6+u4rBQ/w916gCOeg
YxR3kDZl7hp95VDdXMCnQBu3QQ4V0tUVyMHHYiySwpJVFAXXNXN8nDLsRjClsvF+
C8NFdDPbjq00SATLaLu6Nj+E4PjDxPcFIpCIpVTwkJAKU3yMQeb0/pzAroFiAQj0
BAJ3/nMbwYI8FB4a/hLc1eazhmD3iKYKnrGvuLu8UfzTG3GhrCDnhQVwg0XSuvGP
CTmvUeLU0efPbalf+ebaYDn5b4jdQ5bWGmRNdqYME7pFl6y5uewEWyWiKxkRVFV0
TuoBTHXxMZ3cwTVpTDh5ErqwjMEtVktCm2UgiPhrGCXwbm/OaSLFdOMgUb0WSS1+
jMS0hb2nDlo79/sIEvSUxsJ7LBOGzvtcl44SFptXu2wo9WiyDKTLU3eObjuIVPlm
RNYAqdEeeYyJqEIBIGt+7AcnRVZm73TM09I+J4ex8f9LdXZYUTVwaEnWwp+Psdfn
4VuXcvhP0Noe/RZS+W9Vi/wV48EF6C39LtHJDTruOJBWc8UHoWdvcPV4NFjM//vA
cF0xSK6ePsC4rxecIks6DWCnrnn7aOrVXGKKD/8oxXs/e9k4UiMXHw9fhGOY0i8N
LuBwbIPt5IkPsJl0VOdzdQCtKv8DTQbaXnOESllaDH9F58mW3KQvfPgW8X5/uDh3
wen50X0sIip2tSqvlzujOfih485VrGCdp2giqJODFN30SxxZKJPTwQuqZVReTV6O
hi2/+1l3TuV7lgUW8K8XjUR8O000gRVd3ltojpyyeyhiYk3Si3tgXnZOsrEFiDNt
VrKL3D263b7PySa8+2eGxVO3UyAoPKxmleTGal2pFDo2cU9GnJ70NQDJZvDCC0Qo
U77b+7/TIDyjrY/yHZS9nEQleIez2I5hgOX5e4BGrbkzpJH/kAEKOdPy1M+HAITH
v6MfvKOMRKqTzqobclTXtQOv0bc/SuXelNISlixWgtbWzJpofNtx22EFyjGChEfG
0ZuJyNEHInF99KHpWqgDASqTc7WJwQNNQx85RAMXpR0oKxA8sTwPHLipbfniIUXZ
MO5pHZPA8WZoyaa7uulunkxMsjwA9kSZHDZHYlv1MPtUe7pM7giBYRa24ygQTRWZ
VMgFXZmuZq0FI+FOHAxkWh66B12XudGdQYOJR4Izb0EV5pAXkVEwL2b2UeP0IW9J
h2HFD7OtSathv7/It1Od0ZWNsw8HumK1ThLFQ5IapGjx/oMpaQaggP0qaNWUDG78
KVG4jBR0Epz1V2aTAe7/Ecc5egS8apkB6ErDpTuddxzQxNDyI/dXI7FrbEi2ML93
wU+abHZde0acr3SdFdKgqz3ZF2NxaTD63T3S+YahdGF3raTn0KgCJxOoHePQYONi
iBp1S/Wc/nlFc+ne5A/p5r1/+v26yqgWdksw1Hkkw73fYY5lAP7CHxS9cIOBTxT+
EDA0HuBKQk6WFrCIsaualjiyFNDlPqFlHSQ4aMm4NcFZPtiW5b65Gp5pllVI1/g+
Rnff/4Oee095kioUEhpCw5RVk+toYzAsXv3CRI4relw9P0+lnqveau2G+vcQVH7D
AN+vXKDZoqxbLnabyEsSKTtmC5a5VXr0lz6+hqZl5yK7CDQuM509A3yigttOlGZF
lUgCvBDeqzS27Wc2szNrbP/jY7GImHNcIbgFu6FhWoHJ0/mhJMNbc4FGCx9N4jkR
8Ade7M1yWeQo5WIKc1df9IWexMtp+V7t0v1SArljohlIyaaOshol67goxenzaoii
c8QXqc2vFKtl2G5uaG/XAKQ8Wk91AYkELI3QZyCkXkYuydke9lSaBO4nU9uT7c2N
ol0D+vowUFbV2Vzi4eXWQAbu3NObK38OfQRinIQnIL+pmVDa0SsnzhgFDvyo90mK
RWEQarruzahXYXxr4lw66nSP35yp/LZ24vN6hm/XMtKPwuo2m6YIKHe1fiTlccbG
KjUc1KCd7TTG5MpkzoOqAQiEqev4PVktsGEYX0oLvjYdfKO3Cgd4pj9vb9+y8D31
PXQpPo3aFeL43HyieFCah6c2j7gM95UqIdO84y+xmJbvBFmGj5p1o822Pc70Gm3k
P3evtGcwLw49Nk8dBTs7KElCPjtRLjwZ8SHP2p7Hwn3EMxn/DngDz5yw1grHTWHO
Ao+g1HgzS6ERXJP/cKOpru2deFoOTpDsHG8ZqdS36ERP4N22Xzwqj1Q6hN0OcDr3
w4oWUK4PBhZ50pV1/f/NI7twclJvSRVsjjIdQyor2jt5TSviD+tQI1arauoJIjm8
ehmTTE8wYXUCEKfr1nelgZXvIE+1dIchJRpsqi+JH9JmsCQOHUX26p8Dab49c62T
QD3oQeJEwPJ+YKs8LOrYOSDb003BMQH/0v04GuuLKf/aC1lL4aEoWLmPS2k3M33y
hM3uvGvy6dIfs+SoOfUqnlz/6XvSy4DQzeagXgVLdizv6MAnyt6F9bphtNbnNkNh
WrvmCsr2iCHwqbE4LgxecWKM9FXiXgGx19nhdU+agzLPnbYKnb3fH2nwxmhQYSVq
ehMFJlqGhsmhB7NT/uCiIEpaGIh01YkDp1CvroWlMSdZS802EPPXOlIH7ATbxfa/
aEf9ke3Y3aKXoYYAgRvr+vTjxLSAXGdgK3HKWBqWTkKqXdKQQ6x27MHzPKYADL7R
DJrHuuIq6bR5NTVzyYvt893riBMFhutmzkzoDljprUMVxudR34hwWzAPcxoIkSbZ
dAsnPPD0K2qK+kozpQ1s3L75A4g5GADRi3bldfppxVB001aIYPyBRGmk4jDOzii8
m5MnNHWvyBvN8I472s8VhaTV9FCjeMgvIiP56S6XRrdT75NHni3qHc2fM6LE7xpV
6GCcsOojO9qAxqf7RoJnwXAtXIuavnGyFheld7nNtO6Z4PPtbv2SbSdmcI9qKHUC
3SqsczE6yliuF/jW/MWFm+nt3Cfhf7G0XnLYyFHdIeyMBjVXxc3PR2rCZkS/c9rP
uKqWs9osVZWSKYe66A39x2LzDJedLviEYCe+0/yYhTg+/E5G38g6zzMQzd2xWNyM
z+IXo9Iux2Dncho6Lj06S7Af9oHCQMl9vRQH6+/LTrh/VTTXv+UVR7It61+WufxL
GEVvEhptDfKFmwYBNwjrBU+wr3uQXwrlHlXn9tDUDj2lRs8E5YFoKrC9YhfEXU1e
heVAj6LEhEzT3nvU+7f3aS0Gt8GLbcvWon0aEVmkO3OaJSbN2i2+wqJYL7Rg1EzL
Ij1Pmayq9lDU5ZKgnL8ZTvaWgupSXYDOnq3ufrfGl8ycbi9rDz/HIl1fMyBlsrco
579u0yxEG4Ey2TCopGhsaA2jpnhDs0MmurqKaxTfbx4lZZcd8uDzz8+euisLl0Z1
fD9+uqY6mw6jALWXAD6J4SBGuY26xqxmAmmVAga1YjTOn2iVn/kFctlDWJKipovd
WeSwOArQIumDh8R9MmktggWRIWiUCeScr6Z0GSuh+NlARrT5k6Y5marOqilH5V5/
SLqjsa25+MnAKL/gu0EWRfmE3Zux8jXuD81Oagspc8BlN5pqNPjXG2Ho9cbAwH63
n6RMx2ShkC9sQE8G0LFr9+ybf5hMmNsLwjttPAMgL1PJzP5aIlRYEsT0mWgI5dsH
R2XEQWKFKh0hjYGhKqT9NSbCV7+lN9/popgc8XRLcLjnHgLGT/K93N5qxggXDgyb
pd70JyD+ecWeCUR4q6HXVlN/TZvjoMHwCFjXPLeA6bBnbL1X1lqFsPWjyTnKo2aB
yquNHsIfWV/BEl58b1SR2Y79KTHWPHgvm+GeGmFbl+y0R5JeozLE6JJ2DqjEWl2j
g0e+B6cxpD4XJW9bDwPHdbQnnUmR2rqozSEdRpAwgVzYKh9u3PKnsq0KdyBCq1F9
gMy36YguENv5MWC3CGyblDrUVrCWMhYo0fNlYky1UB5uFpyw9RoIGIVZfaY5ycR+
fPWYErToW/hTp2vvvJNiEXNobIEmMJhcVpA6Nf6uyOIqz6hGa7AokuDWa6JdBbwS
uo3VJbLh07EGejFXPtKAPfyFT5iirzNwnwp3kKGzom9z8G/iheq6guZznCcI/91x
SZ7YmAqrkhwk9F5tbWOcnwG8T2WQ7vejXmUQwexEs1AVXujjuuwScbY9wAoTmMrz
ktjEy5d08RWN7Ehw588IiLkIzrB3dSte8mA6JVwMqGekFh6vt5ETByv34JfrwlnJ
Sht3+3lPMxrMfbJqHeKi/3c95kdf+t5D7cYi7TRd5CemGHrHmzWWvrBDbetG1aaW
Hjskdsj8C1obFy1FeleUGd43d4LIp24vpRYR6wSciaoDKhP1gnWFY4LJp9D21kp7
UNsJ+CuJuB6nITYeRL+/IS2U6xoJdc/GXCgcgKML1fOKmkYbnxZxpN5hf4NSP3LQ
4DP4r52l2kqUzOCwcVbhLVRdnaiS1olvFHu9oSjXEsRsepPybJu6b28viy9Zo8bC
glTWaFnTqxhKnJIZ/ZBUCVI0Ev/PotwsR+VqHP4LT5EZdRizHdueNlw44nPog05V
lTntXmtjC4iDN8o8nsB2OLhmKtLjg+KdewyblFeku5c8dO/zXW4LJm05TsGg4YyF
82EAzuFr7yuTWOyFjcz0Ilp/CTrR9DJi6HmsufyMkt/n//vDWumYwBO9+yS4Weyk
Lgn7YLQ3Bqo4UQoDaJJAsAbq2eUHgQAZ6dEMoIeiUAvEfVgMWXQluD1iw5/g9q73
rsYWqD4VmIhtcp+6W7EmRXCgTM73YJhXDMuLUJCOTRw/t/0rBlLS7xdVRbop0+iL
UaCMAaEmdxHwychEO7ZwtxlvS42kLdeTQQanY5lXCGT0jQ6VzXN921lVi9u/NezU
0trNN1Qt5UPr0lcmReFZzv6vn1ksX/OwnQ+a4EZGOIG94eo+rfHyysom/8ggkQZE
m9jSIrvx2QQ09k7MzKLUBkHVr3ZgsOizwxYJfO7eUqniRwoFSxvFcjNeTb94/AIR
upPenurtsBfjoYJFS2BTITdZShY0yd3niJg95hKNouxAk+8krZSkQ3CZjWF/dUOl
IgleUDJ/8jGwwAHbrWZyu1R2CZ14REuCcItQNFSSqjK8gzcCy36FQgSXr25SSekI
KCGbGhIpPfwY9wrCzueuOqWAxygEgS7/yGg01eGmMqQ11iktuDogIAoEvxEFcgTE
fgIcLYgswDucOiKMXjGlhURJZJpb/LXEeyZTeind9Ma9Zn/mCnTM+ltTzm9H3joV
jUvKsC804U6e1vE0VD9OqHHVdb57qjxmzDRteQmaKeLcOLqj8RB0t629U0TUgDor
gJIpiK0If4Ol5HbzDVTdbva8cU7ESgngy8hoR/JM4HAX/8s7i721Vt2lX9ZzRQNU
6SLtFyJ0xucCENBes8jf77WP59yyhsCQynQ0zuPJbnVx6Y8dBuOnOs7rxlGYQt4u
8FbgTCoKRnJdmnRvUgzFCOoUFRgqLB8S3+EMlqlsGa8DQLkRaJ14yetc5FWxoMYA
tDQ/ooYyOpjBRDjlFBGxJq0v86fb6zkg4Q7coSsIgh9X857c4ns0ikhQHR9LZGMq
1Pv/GrEayqBeSuKE3GzLQAYMOYTD2JGRuz/fLFeHIIa2aNoqH+X+Pvuekov4NJhd
Ayk5cRlPtnteWZmnV5g85ugtWXKB2+ZjiA0+yvWz3+rnnda7xqU7KCXzWHWj1ihc
9gXVPkj4nLhDdcx9VagZEPE/i8QprOl+vyL9ubdGRE6+vdUpCgFfY76gZ8D8Tkf3
rRHcqausmqk9pAoHx1l1iZ8zCnvOXw38vqqX32uvBe3+WjKJ4stlNqxcp8aeexEe
ywl3AUO/j7MDgPB4q89q0cbez1Y4X4JodvNyRo0rTOziQEbB+fTXYUfbM2NX29e5
jO+FwFEjtHoe637gmTHNeIiyapG3NFpl2YBnfszqlcfXP2toPWzZrT+fU81VlhrQ
/HSkOAyeGTZd/vS4X+S66CkrN/EaLk89KxyjbkrUhE+lTxMv5UcI9QcZAgRkSDXC
5irAJOrmqibxrvwWEpAzHzBimm1ecLt6isyDKqAYgtAPWDna8qk7l9hemTOePlmc
acebSZAv8BnYsYTiQuMD9vsTqZVzfjT9eVhuYjyOVtA09gSCYrcUuJkBGhMjXzJJ
EhcE4+/kMIrXy/Rou2MA4bCNP9fOMnERXdiQarHypyiYjplsyGPcxeFyYMH1n4QG
PMs9qtZmm51j4/mBNf8IIS87nzzkR96IXx+m7tLKD3sgfs6uOBeM47PG0RLHWIRh
TBkTHzwpZRppHH7aC9RD2iuh3jk5WsR+1GRucgm7aIFx/jWs5idfXGiWf9FZgkrk
GU5OllB2rBjEzgoeK7gUl/kn3QHurHWYZuVLkoGFJ4JF8MzxFqSYXOQSU2YrfSen
7qWKCAAirGsC+c8AoUaLZG96OKqD/8P9DK1a5DQjT4efXu7IY2SycjRsHLmry3J6
LQewvzozagZULSVJQ4gj0X3tS9diQjUE+MQ27/fxrFhqwDcpLOWddo3G+CfSr/ji
KyMXa6EfPXNV7OzUjKcjvydwYxklyTp/Wj2PsfscOEyvKqyU70HfgmY7b5xNhFD6
49GW0B8LyUz/g+KDTSm6aeTOgQj9BNy87EKmHHBLKexYB8l4LAGCjsJhhf0MP7GG
EPsUyohDkKlQy+npsMc0EpxtpwJGZIbtatQg4BQDOizn3lqRXbC+2GDkAKjJAWpe
CdgpoCHbuArbstey9JXLVUu2DUBooDtOxyjFKg+koccTN86IhUkXAdFjs5ty6ayg
TB5h9pawxb5zz8Dbfn3OEiTmClT5bqFaAjeXo6vjEjBwfYLUasrl/DGaUPiGM5fZ
OkPkxSJveSxS1wEXQ1hpIK62vS+m3S4ftQSF2jnreWbY77gZIPmREFhr8SLzL1om
ICDmXoTG0DJZGUKbUYcRPOqc/ZZR9BKLzfWAwRAFwQ5GCthmXls7BHyoABnMIp5R
UfNUPu8f8okpBwE9G2FMpHdsbQrKf+np9EXRhc32BXrWgZTZFY85794ZSGOf9Gow
a4scBQoQwMjWVkEbWTUsYM9kWJSeJp8XHEr1xA+YyF3iJZqiGyQ3nSZvyS8SwjcG
9QPGlEy9fR8KGkZlsY+jbJVXfPqS3ymCc4zVpUYSu8JKeALkJu2NonBbwP2EvVvr
zSL5lqE9X35RAq4vrEJMa8odmdLxG6LYX7D4A1HIIP7bwKvA22Wj1U8Mz8+QJK1d
TXhyu7uxpPgozr1GfZOF4wgQ7dtFfHS7bp90DCqktGo3B8WHQx92u2+gDfOk//We
F7DpnP9ilkTvi+dylKqsfeIFStRHYD56CDSgI84ApBNV8RXHpGUXmde/W0a7Anrc
Mzg+qVFDGvh4oUKq6cs9bJn/I+AA2c3eIjGs83uddtE/FE5jGg+SSMYQoSSgFkCD
OTz/Ize1nA2VGotcbrN/nvXau1b9g99hMR6pBZ01RlU9n/+1cOTGk9ObdDdrwOYV
U1NR8z8WbYQsqVKJYt7CFisM8osVqZhKqzBQ4qlRkYPDw/0Fq+1vY9lQHFw4R+C7
062R5uN1Bx+pEFAIs9ybjqEuUGdwoFUvblwjNDzFb0le0hTHZpPuJPJLWPZrAD1f
TdIlzloCvZCN+IpJzIbARhk9z2j11w9TFRw+A+go7RlG5ai2I77Kz4SxHfIXJ/Mf
q7DoLR+/hUjZ3y0Gm9cKBxxm72yv/CZW/7xUPIqHc/Cy6vDFlKftHMKz0pV4Zk/d
5+1Ms854W60nfL5QhHViX+0gGd5NWZQPi3b99k0zGyoVzAo8s71xc/9zZ5UY4psa
17DStwGV5z5abyevfQldZrZNImSyLiQycJg8ulDaKunZyYDOuxpi4z9jfLYLQxAm
APoeDiKs4dRb9Zm8Ts/Cj64G2f0eIENCpIqhtj2D3BSs+IPDZ5KyLhafUDaVVvNa
MBz5KZvQq5TiSwkbJeY7SftMbctg1I3RJpKwR3h86bjvT3zbjz/4cLxd/9Q7HKgR
wjTnu/SwNpTBfGvVJTwuV3z1eR84GaFvSnmjl5e8kTgnPSM/kGtFOpyEArsgggDf
JMx0rqD5boXzaL7rd6X/98bOorTvfWaeLP/pdr+0Dxml+stMBCK2DUx1XDfkdNgV
72G8H90rj0SrjOOGgh9j1q0c2csNuepRqWNfOFt0T6zqR9Mvykj4f8TKXHMeKH4W
crx6futEvRwEDK7IxkZtK9KVzqHAHhZihN7x9gTMmZODWj//9zVz1lHXTYhOguNv
yLsYu3sk2JdJZ0EKCIiavSvKPuHx0NlT0zupTjVtD1WCvAPzHMUXIpJg3P1hk5v4
hb+wuswJihnVoGconV8EqEzbVU/8NGOoEYqhMlMzKe/+YOMVdzgtJ/vDcKa9CmBB
E2UpN7RBoWoiahTuqD7uBzHpNiku0y++DVcyCSmpYEubMATkxoc4f/jdmPrgrdHG
r5pFj2qWWA7SeUNClVHOIHl5LRkiD3LfQzGQI026PuMANft+7JBFFGqtBogzGx7G
TCN8BqHY1w+WEBOEEnDS7dk7u9maxXL758Di8tuHK7uKNhovqijGStVL32JIg8i5
K8m+Yo3Da0m/ZwXMRyanV8+zKTMySYqaFsZMa096kua0reCpRoFCwgwelCtdm0fD
TBFCiggkXPYJKgqSuTZe0mw8o9PKN1UmNgZzi5aLWVKwGEKU8nHewNF1tPHV4aEY
Gm+wND+Benib5rUf5DEjJTbz0E32U2SQFcDBzTrtVkJY65j2zxCl7nMMWPHZEk7v
PHy5dc40rDHwYATh+HjKl6dKY7Su1aguki10mBFQC2DUG2zOtsbkvYTq6LtTpL7P
MdMgjh07enBo00K6X3a1kS13hBMM4qYaSOyVctdJ+gev//5dJX+Nx38TmH3hiVYk
/SrAHaChvpxBfqy8f4G/3YbHtBrNe1ri7OloDDUW/nHapRHte+YGjpwd2ADCoIyF
D/uGd1roUnZsXBpw2oTPdZsZVPUUlmwDGDoNRtmJXPLKL8/Kkak6YDs6gO2YE+P1
giABzUJt2lXruBnwJ743mfvQk8E6pI2VPUd3AFrdqh4DMalfFiNnAVimthNUoRVi
BC5V9rj2azuPVu8nMXlh5Di7PFpnR0lsfrVFaGcrJcZhNAKqtZARru+apI1wU1n3
rmS7+7kwQvZ4UhvX7Jq93atFFhG6kYBpA0/fmbpobm65/3KTZKZL3JWXQSE8Mjct
BWeygrqEWfyjpNLWDtG2kfAY/r/G9mDe1pFt4VeruGT/rasNVVkRAe5pXO446FMk
l/fBAGPliIFct0i8utnTCMl54F6NVjN5hLzxLThMzc/UW7RlkVRTFwVxqK9zuH+f
InwV8lyuWdnbpL1NUOp6Gvh/hnHYAciXpx0D9Bc2VvQbjI0Z6f/GEkoNKOxCh9wA
JIc03NUvHPfFnubQt0K6FBf36yaiRVUSbsrukLbKQCt7SI9Y5wt2tzUmX3DUurCS
uDEvEtAo8/lla3cwKjN6LZY7wfhauaOFhFEtwnu4UC+C/vcNbAonTbyziaX8qrBP
8K9sZcveybmqMUfzppW4Qy8z36pR/wvZZ/VOwoFnTWy5x8T+vBp+ZvPbV6shQ2Kf
gpd48WKriaKGOBicjRggLrmtG7NuxX/FU7Qp6sJkylIzTFWMFfBPg51rmBhSajun
U4U2gmQbV4YsaUKAtBRCSIu5sxhT1rcWigEpqT5PXfQdawJVpJmdHSMLFmqIOUfm
/3/MQaUR9bTgRk0PTwdCKeDGPtmPF00Oy30Ch3hXP1lq7E38XINaCSgagLmtf555
YXXdRA3PC2OTML12jmfowyyT+y3XNHPeMiK37wKQoKCbJhrGjboN3HniZ4UMG4Zg
FJoaRm3wNQfxo3zOSZSDth82/3nmTHujfhE9OcSJXw4ZomqnCnk8Pc2TcT0aQtvu
McF7vSqT2SFowu+b1UHuQTI0jXz4lrVfMShbUFCm8UkiPqje1MQ/H62kU6uVfPXz
sS+MC0s4cyXYTzqSbtTet4LYtbXH41sKcEwiobESasQHAxlAWmmVmNijyJ3T/WiB
LqFRMsyhGLY6q2L0rm9q9/DGuWKXVFzTefTcJ+mSrshO25CnIv5Bg/5WI7Z6ORQ1
snKr4mnABBKBKstydxFwJ85/So0aDV8FWNIf7dlQjKl2Et1WkFzz09nzW6T7D2cV
WCZugrXWfjcI8kpYFO2ZpGmCghc3Zzz+RKJYyLa0ATjgdkVpDMqQop0J2QPr33PY
ts245RUiIIxHzlLeUzgHB7KPO0GI9MKt5kqO7SdOqU0/M3qwVpwHoPGbplCBjkFj
vVeJ4nbiSkfkFu5V+kPnn8KoiotE0DnTi7de0MTW4sbeI1VTfNgrdQVDcPyYxlxu
7QYMDlx7VWyLRePLsguOWt8MMxOrHI69ZrzTalkAKVrnIyfuTQva3aOmpmGF0QO4
l1s7vqWS2sepiAkW3e2YjXcScifV70L6uvFeZPe1KDHvBkA2il9AdeNHLaJD42mO
azbpKPPVY0drkaoTgFBjgwGFWJz0ZI943YMYQqV6z0ZaDIFAFcx6sOLOpjs+hsyr
TNJtrQRMO+ZZ1zEIbKUURX1z1oNPTmKIs10BQDumi1WzuxcsOv+9IOKgs1ocYWxM
Yz6sUzLPYpKBpyshN/7/AR3nxaucgM/JBxMAflBgHzRc/RxTbtDbr6VioGr67z24
3YCzJxiFo0w7xsl2hs3oqH2dvgngL7W5O7TjNrGKYEziuq1d38vzZNyuM9yxSPpI
8oyENT+5ArEdMSOt0r+vrBcCNUUUSBoT3P81nm6yDnUQ7faRQziYN5ZFa1ayt0Kq
sRM/6+x1NMGKdDbil2N819sWIHzanPu7/Xd0TR678q7F8INjdjaXBZCRAl5hD80s
v7+AhAy4+dL1uQeH0FGHuID6Ba9H56Vw6f9VwZbPVcWSwv+N0nDS27+/33eSTLs7
qvw8EEOE/+r3q+jPd/QrSLujKJWqdilM99Wi4yMU2lLpBW2oNB98TN4cXxrKENIx
zTYKoOtbFP8Adjo9934XO0LiGXsF7lA01rvg7vukbAq0tGlFY5dUStDvkS2Mznea
J4glO4+Ad1uCRjVaHjH+B40ncE8GnPTvDtWNsxIGmvz/ccMYj1KX1jo0Ffco2nQx
5mUvQVChQBkREWCPD5f8QLEotA4D70P5wjYRa9MAVKiH0hNcAQwBSEAPIVX9sCDN
L9nprT8UIi0/bVnFt/V48MvIaKZjrpDPoyo/zYD3yX02W7wrKGEGhqfiKRknTzF5
sESd4yJ4PEDNAAbM6qpgksMghrBxj0R+NXWd00jx5xOQU+rQ6qzCS/6t74DI5a3z
zgVljTrJqQgZczQJoYXn0hr9AkSRxVxzQ78udt4Nab+bRsQ9q8HQi/+qwR3crixv
yMdT/HW/etpzuESHxWv/c93/9kE5EkP2mddLy6sf6pPRUZZZrDChmDjs3GOkPdBF
woVT2oyEiy67zoXzCS4Ksk2N+2kv2J036Xyx7fimLQ/404v5QYVfIThFeQzSvyIc
J5xn7bKJJbprsv3BU86NGJ4RxIDXV9cIuDCbMPX04kKqdhLPIyS+WmwJJst/i3PA
GVQzabybFfLol7xCfohvApOtpW7+nw0Zicgpw8PgJax7XcfQKy0uY00JcAlEo2Bv
UEGPU/2x9kAoR/DKtlTZjtVHHKt+Ay3AM6lX3h1YDDFfLk3Rm6ut9iE8Ba2a04T/
blj9VS2sd2nhw3w9mD2JlYd5PmgMKdZLSZ2K8Z1gGluuReOdgTojPhmXi66yW6PH
9nRfmrvL2albrBOnMIYr/dDG35DSiz1j+9Aej5t1VR8jKFaN/zpJt+1NXFZ/Oe0p
n6nuWUwG8jWc7XrFd2qhXbvg5j5UTcKSbRI3Q7nFbIi8JeDti04fw00NC+OaJ1nx
o6kGnSr9w+E95uN2oMR0SkqRJIlgE7LCKUMlVLEsLJtCa2ElCSyNE9ih0mNWQL3W
nflzC4QTnbDS5zdVGqfw1HBTpNCAgCgu3QdEerdRkgYV1+ZQ3jRMojS2iziqTg6N
OG+9OE8R2KY/0yQoVU5r8glo9uulIWx0NkQnMWG61t9eBpl3/6kwUy99odPKnnPg
wAofZR0otTqUJ37QTRNNWYJrfyn7l1LuDqvtY/TQokMqqoICju5uWP6zG3DV6GOU
/RQGR7J7wsxFjgeJrucFRZm05z5KcLyjmYne/ML8oYZrNxWPGvkOngvo4QsLJYfx
dUpgOMwjrz6h74hCEIrsDnkC6wQMJrDWvsjXOcJRy4Dm3BrzJ6fsLGUWU2dzMWVq
GlJi6UV9jtqhHHj1WZ/98eu6fpAknwVMfqmI8vxq7jz9q6K9fRaTzhiEus9p3BY3
f8gchjjZRwCmA59CZ95B+s/piOWfPokYfPMYVtDyzYgNkF6H3RrfkEu+31pvLaXO
rdI7mTeeFVF7PInvE7Bt6J2gaKFQnaSYfA7MAO0NRkTAm9+1Sobz2KrpLyTTRejG
gJyY5LyJjsWSb7YPK7VRd+K1VhN9a3VV9LQKMGo21mmr5vkuPLl1gXGtH2uwNxv+
qrxxP96MMNNDZSTgGeT0IeSpI3/8i7816gH2Pj6FPyIAtVX4WKR8J+M/hQo3/bo3
Rhx+w0Rx42U5rWENQ2pGAAugBKwoCkufEGk0TJYUx0OJRIP6gO2qLlsHxyfnh7MN
9fM82HKRypugcXyPKwpJFX62VWs64Dt5WQWN8NQcL30OOklHx3EIXNu76q8cHjHZ
1B7PVhaCoKL3XcTMVWHfGaZzr9kFtm37+ViJ1Hrb+6Raoc9IbM1r4LWRZUFqKBfp
c319vR84jaLEBev51jUGKop1CrPeYTnpCBXG0IGFopiSSUBfyledV0+sa2iZmzWH
oIrktD2BwERrwZjenpCUbkAkqm08/nZEm2FMFKxv02ZyXG8w64CBJO4UD6Ugc5Pn
IlB9F0cfH//HtWESYB4dqnMm8zJl7lp3IJt+Z7rQaKU1ZI4urr/sMnVsEQIMjzPa
f11atIeROLSeLghc7wrrXRw5gPi1ZZc2BQKH3oEccexmu0DDo8wR4uUIDlvCXCDy
n9di9FD4RpEaqL6h5zmxOkMg9nLm2oaympLcraajMrjiDQklYRMZQCHOiR45Yuk+
beJHwSbglA+e1OuUFBpIcz8kPdqBkCe3DhFwACIQ/KxnxjG661R1ePCDXcLdIJfC
UE79QOPPoKYnX7yDuvLYj92WcYXyjMIR6D9Isjw2oO7uy938ZgWcXHyiB2r1Tzib
EFoYvhHStvz/WUSmQyT49V5N1MlGIqerr4nRKP6OUmN2P56xtXsOjmwhfMA+kVsy
Py25jzc19XsnJ9uR0vekqStx8LTj32Y7AbUau1bjaS1eZRS/Z8Mm/oh5cZzyAvn9
w2QWS04VWQBWJwAqOdwmq2cIYPlXA4RiWggwmiND2rejRrwmNFWHcp8ZA8klJRfR
cU0aKcoINOhKvn+su3WaouCwE5EeHTYXP4v7YxWRo62XXhukmPYzFsUKsns16/hy
i0ahzcX1d1UJh/45H9BwVqqJ3cFLfcf7G5cghNvWu9gc6a5LcLqSAR0uTayoZma+
aG03rcIkDr46uNAmldk6rBTd/lxxb/xnmBbNNCocxwgecIOnu6d4eIzWUGr8hRPo
8UvOQ37cJJMSICMzBZGIBfd4JTMcbnIwWPR3KzijJgC88fsVTYrXi08+ne7MoxR+
a24FzA72RRbhRYLZahl9NY7dSznj5dbYpZCwrDdsMBzSFTmarYCWYldDSKlNTzRT
YI9cdGIR5qBxK0+JuQv2f40o/GxZKpjyVeXf/9V4Wu8L7XcAX/SeCe7SsGYTVQ6L
IoCzDwbtZXJfe/nhCUtQUeOvheGRmkF08SckCOh0lThWob8CFIOQjBwV7YEn1u+u
cGvaA4pnSvAsgrvjOCj28vlNsNakex/HEf2FYQAnsck8kAeWg4ZiB12iReMBn38K
DGrIHd360WkgbnWBWmpDnebMlNoKvmRriDzGpppiWGcbcAJpWa+A8mff2Vt2oqnE
5lWYZXwu86UXT/RU4ypmoZPn33rHmGaM4h9EWxq976trvcB+rLqmGhlE/ns0UaHg
62lsbNUtb5LVIFs0GtVnz7n0tF9VcbX1N3IMLLCaeimxBfZo2z8YnO0CMT8Ax0io
Amxj7zzElGqOkqvgoxsvTUyBbARjB/W5UsLwCewk9aYzZO+aG205K91edpJhWWue
m1Ol9fNT6j8vfkWCQIqsEkTEiVD5InPyQ5DlqnAw2oV4nKXiu38W78F0rb3/5Vyd
+G+yrw8bONciTM7/T2F4DSme8icTprgtYIMOBddkIA60uwy0RDfok+Z0OoG7wf2n
bHZY9XWwUwIfHRRj67jBOwTlwoxG2tS8H+QRNoVYtor36GkDn5djdCNLC8mD66aa
vauVc2sOxO6wpxnXi6KbvX46osotHOFcAdtdEtvoL7mFEGIvCpIqrpudcq2OHvya
zFG72UynCbWRdHrltBVXRg3BXPqnVIVeVFuhGbJtRV90/0yM7i/EBuXbVRtR08vo
bfe2BFa5Zmthj3hC9HbzxvR04y9P6CpjmYzo9PH+no0eCVFpA5Pqtlt8nT+6rvOq
4eES0TK6Tb8mTIzmoDmmXP1y8pytQE14cnFc5Pu3xEbNnYKAgRxYpJ8ZrP7eJzXQ
OxGhlKW2tX1EKtZgkwLPHPZR1UBfQAV73J5CnIipfDVotLDi1OA2uddjvgqSZaTs
+mmeAl8djAYB3MsehGQLS9mzBlDFMnm/w5sh2sv4ncquVjrrDHzhX/jk0pbv1/Mg
p1RiCr/CiH0aXSiMWdIFiByKeqmRGhrF2HAMF4T5GFxBIj1WIdSgNxbmLPe7xscr
iGEW2iN/yUnsyKNImmEMQBNLfCgmXITU6TZQurTbVmu9fKuKKi5tTy5SEwvs+R8r
ZE73VQ4If9sYiX2ME5CWeLv5sF7zWGJZmU8pvMMgTJZgvbnq2M3MR7IVNWJzX4vT
TLBrGHnbIdOBMBCTAW9DVKyMTGnNLHGmYJZ7HLGpRpqBuc6iH+c65RrSKQDcz9CD
XsALevVLIANYPRLT3g/s3l96id+X1JbrvjffESo/H+szbsNHKf0DyaptOWPIz49O
v8vUqLMzQWXIMjf8DTAchGXclKi4Rl73JJatbNHr+YGoClo4tvSBDf/5yqUUad8z
lljFi0wN7RIo7uSBp+QQjuTHlL+rB21ObXQHcSGi3Ixv7eU73OnQmzeMCr3Ug8+v
ss9qyt7s+dEjG7OIHamN6iOK/9WvsLZE0rHB53sgSYN+31KWvfV8LSoFN/2CsC8Z
YOdI4OKY/XmEbh4ysD4i/wdXIUxITyAfpXFVwj1jNvnIkVPFZNR+ZFMvL018g3T7
JJvrUGyKfUOg/q31viIo3j5O696yJGIS53OCIGB0Rlq5Gaa4O0uaps5fl3yKGxj4
/MeB2rnOsIvkUwjR7LYlzjSBb/us9z7W7iordnR4lKDJgpw0fPsKgjckEQNgNKxz
cqoljFUtcvK3fIJHkekwA7xiNO132SU+/q1deHY7isGVNgo+xasPWDi5soMj87Mw
gvd3BeCMkVqtQpqAQiugLck2G2+hhAbNQZcroVVuiMcZgRGOYgo7D22svtSEdb71
FLC70oOlbsucX02jGC9gCzskO7WGqHgYfty9qUkIAva7qdA0ScFGf8pTgFVBCXEb
YfmSJZJptNSYYmyUGpRhmLp+AL5BAwfvHGFwyOYaWpturzxR3HQD/sVbACUnVDsi
LEhgihMZkdBOJ6xT5ljMOVQTdTw+rcwuDnHlz0oyCq0r4wCbJT3M8JEKxlkCvJ90
VwfensomRjoGVONBH2ansYLRusLdPOOBA58NGWZY20NQ6lbxemuy8LBtmVbL/Q7O
RWtKDgLyPtNpDnvXcy+zSPpy7Qp/x9jE0YzGZVCzuAhT6hBPP1SSCEDL2X/CU1j0
bc9WwCX8IfZ11i2FVxx9OocOheUzXiCPhT0NJQOFNrpj9roTSlIdjVs46QKz1hcX
wLvmwlL0DSwqbJmEuheps9M4uXIEwhPmypFgpyqqYmv4S4gYbXLHM2+g++PAPeoA
4XxYAf2M2AtAZ3LgdjprxgXw+yunL8NJEm1xtaHRtrBWhrYGbIpkpucmKuZBLhBa
aSpGsKgHmHuYff4jM3gR6bbipE99SrfZL+eEs/Nw8jf+dWBMsGgsHClTU4VBeArN
Wv/JqFWrwUgoPJVV3DPwD6MWAvmPfj9U9CrbnXOHyfTEwDPVXJAjRo42K9nD45Fj
cSd0iwh50Jx65IJpLC6df3FnCzKgs5SvBqStDO3x06EJylNmYuodWO9sYNME3GrY
zPmXk5w9JQUnFLjU4NXK0lZWpCR93HfBjiw/F9OFAHzphkTM2XRQUngDeC2Ms0tN
TKKeABig+AjYuT1oli+0OHMM0MXy1Bq3vJy0oWyFRufJWTs6xzXnEHXNEr12r9jm
rF+30Tt79frfQGxVTSbwgeeZd/Js3uSkhG/6Kb6DS1rIPO9cbTGd/+oq1+D22ac6
Bwzolm17CyKHQd9dm2UM9GjqTL8Fo/DrOqWqf1dCuDV2pVemdsdCP3rzQSdHBuOg
oazXzxepvsI0NIdk9CW/bRUtAKXiqszXS228AfQMK8pOVqYhocfcuT33M/nnz1xY
yWJaBUx6vZabrkv42sZqxzcCwRyWQdQW88YfDti4HTBNlKFg/cEZ6pidM+goPICe
7ok4+09JNC3Jyb6JsXZ+ZUF/YgvjIhueN7VKRTRIv+NL2HSea9lz2mduX7/1pG0Q
KT1S192ZdWrG1k6/1Dm4jq3GkEFtpZJUny7ikcnxLg+Z8f9+DdU/oAkjUmfYnwJQ
pbawryhFSjSaFD3YCbf036ij/wrMIZfqkNR89Y+08xN1bVO4x2jlSYukLbG/LGuF
PV1t4SbgG2m0Q1Rm7NrO5lf73NjziShKTX1mri61V/ITU4q1pgtHTcwtzk/QDqvn
YzsNvi9PSJibRDHqQFLJTny8eeFVnA+aJxiOt9VaLzsCjBtiBkK75qTR/FzhIE7L
XzSHGUFglk3p0MEKbz6NjaWrNR773RRKRkWToJ6Vf3kof54I900LJ2d4rP8W+4xL
Qbtzm0zks9nPyFRvgW5spBIuOxgdboaqF/F2qizTFp43m8pCd5on2EUs7fehVagr
wsgLog1zkAvKOMMen/a8TdY5eDN+Dfax7WJGhX5y6KcFcm2zfeHhaBxKcZqGkayO
cGpG27+SNhI6p8KJID1Uipojz0rdXvdBOEfmeLAdQxV5Qrb7ImGdj809I3F/yMTQ
LmQEpgUFWB7ckh5y8NwxgfKG5nUfLqacod7v00WHQlQZUl8rqFmGypeTNKAqp/dI
kJ1k8mRUlmNABKnpIkd39uVY8b+mQa8jUwgRKwHUpT4/LqKID3aeoi2F9Pp4LoOv
x7xUS31Qr7Pc3X/LOnYh2pmIFFsC2U/tzsyqPGXaDNkbC5uFGEsVtl3HXj5TwQXc
3Nr8tETfRQKJ+kdbIXXDTFvT/y6xjGcX1o2UwSV3p4BY5oHexVwBhMXZzNIDkJS0
IDjtbOV53QCHpLBwlvS0btFJmEg1v+kIUArXJVSBiqwPPtqNwNFPj+tfAXUPjJ6u
EBau6fPfCAUSjvsgZLO8iXn3H4PQox/3Nkf1YKkxM7tgXj3D47HsDmzRA/gfpiYc
l0AsSseY4sm5RWT+OK9q3p7+E3W5CEEYTfo137Ill2yq4TSeUg9/JMHH86GSfW/x
p8Vu+aQSxlfq2jqen3nEsIl1HZxscl+GsL54itnIJfhf0K0zFwNhWd6UZ+Oauhc5
4knc1cXIiK4x1tnfw9mZZVqex1SGgAVQuWwnr6/Rwp9lVzt5kLnGMs91YVRd9Xog
YObgrNx3rpivnuKJLKgJestDa5cyKDKCrrRb5lD5HrNxawVCR2auJ/EAOii0Q1wk
nRRyvpPQlCvcV6qFwp7cInyOjM8YnRsNtrlsbm4wsM34fu/MOXIJuAhl1RuFDQN0
3jHFXYa4piyrMimnX7KWcBdInrwGSyPRITc/Fqw4w3Pq0jbRdcf15nS6kmxtCGzU
sIgXNE6+T/kLgdp7mRNjRsHx/iXbIhLd0JtViAIYXTVk+dg7rPtMPADMb5oNc8Ga
rziT/VrGBylQNN++ppLyNw4W2XuDa7LC5KF++G+EKix3sppd917bwSugBQO6R2Ok
f861Xy64CzyeeJYRbppL3enVqhpDq9iI4/tvl2XoNCchLelP5rZbNVnDRGLkeWh3
TzVdTw0ZY3SQdNq2KMijYXhK8ro0Qpxrn/h0gW2auB6uVBZ+u8k8zK2rbjk4klbq
4qh7OMZkswhM2Q0DYMjbzjbTaMk9syA8wRK+DF7paCkRImIIjHoKgfwxUTHfUXkt
/ghBdxT8xcBx1Uv7FHIm4sXz60xlf7lavT+3Id0RRvtn6/fAeu6bych6M5E/VB8D
PbBezia6J23VJSsMaLmNSxfnz1iCGRExIW/P3Q82Bd9WrWnu/d5JsJS6fu0WpRBx
eXtRMMaXrv2Ao3CVASGN8jHUeAspZVg1CnhOlc8o/f0cQvlttmtHxZmbCKqPJDC6
zPNt6KwF4NczRlNq7oKfUiYHexfdDps+2eAlPHNFqaICxj5lIIE+pfqNZqoe0vyK
+Nwq4SBIRAYhNjYOLiuX26um5nmejXbaqiyLOsEu5ht4YVTHg+UnRKpSrwlXTR+6
LRZse1q7nmz74Ae9NNft6nm8RnPGQOyWNxkk7cEG7NeCy8QjTZSj/YJRyNPYNR28
v/eoZ60BdMb3j1OnP5gfMb0H2RnIgA7ATGJM1PXWJwxzPb5n4eFcxELiRn6MVq6Z
QEscOPw1jnsw1CnKkYUBPrjGX4BF16R4n0fu7jIdgpXBIyby1ISacWgmIm04oMmA
xInFfgaZZbh2PPv5ZX/BEr89blm/k44WKH2vFDnIJFnoMXW0k+C8+Q3JULp8u757
DWqt7SsVQUn5N2QEk3mqJ6kniuG3kyc9DvRHcOss4UBtEO1YY35QvRcL7K4Aq3j5
uHZuNuFcUOyw0RCMf60MFosjlzIstcljdzI0aSrZTojroZzUOhMUPi9wCigJ5/+A
QS9LFDC7sIaPHzz2i6ME5x71ZfbfOwfxUiD+WfuTNr6f+KXW864sSfvjQMY/UPL7
EnKk0prNccQxH3F6v1Q55fWto5Rc4DPFYdiwyvNtIpVMhLqUfIQwrTlQkFHcp1Kz
T+ohcyGWUgW+/CoRYxGjg/IRgqWC8fkUWS2hPLccgAKtRYyC7Me3bMRAraPBqITc
uBN7WRdhc1UyST9IHRShtEm+JzXy7FQttbn5n0Froo+zkyOnALTnljBPX47DKBvy
Zn74PGwnf2cqu5nBzLUNwkqvzG70J6V+D82dOoBulqP5rW8F69tBAaZYF5GKCN8J
MbgGlcaImqzBj6jQTFCN4eTdkWjp0xsdtPiXkp6skcMZJkGn44d2SakPq0Eyk4/4
ShXgv2o0771kCGQ8qUaPeTa3NUyIz33FNBOnLk6R5ReXFVht2sFwNt3PuQ/lyjXv
N+C11RNavS/dUdTavmnjj0K+TE02AmVwn4A0DQgeDPrMO5AkSkjOz9GTsFHk+w8F
VHSwll6vTIBP4I0pMeC4H4wIc45c4z1Zx6YA3pOcdT8GjIMCr2z5V0Q447bztvMC
s7Ilbthw330+nUkboMzibpasw78U3Vx9FCcGG3iHu8aqiEnL1Ipe0HEDZigxiCoL
2372nw10twp5VNlhJmJylM4gZvusJwLZapVKhawKQ1NxwU8afpojTgZhuLF3wyai
wnPWj8yMZJKOzCFRJ8Iaxl8VAOMCBuwFpbBPLoiYm14GKS/u27phme1Wx3SdEgSm
E8Sg3ap/asqveifqk7dwuIPvLtii3L5u5REPF4L1jkCWj0BdZ4046xeKSMNRMqMH
ioGrRGNQZnioQdj/MIX1waqUEZGl4e3F2zZcm9JcigQks53ESsfp/ec+UPvd/31q
MHIeyO9rgjuLNxnPApt4PAbQyaDAGGioUPvzRDtQNaERXgO9wfrO8VvbdiuXMDp3
SauExOeyuK+XrVndE+F5NEcY/OK3V8nh/YCIr7ks04QJKvcwvui/jjeeazVwL85Q
TGf1rb1PkUt8Igygh7KCEMFFid/sxp+TTlvlONMSfl+MIQ4ownK88SFkAYIN0Ud9
cwuZJIB2kvGFNCEUzGFn704DLphfJ9QTRzDR1+klH7BB1Z9HKP7MsKuVP3bF8NHE
JzgerMUIqxYw+mUwus0Rq4NkGda3p/d9ZuxTxTUHOO7OvNztc3OyqI/Ne8aQpFXJ
iKciXG7aHMwlKtGnoNVnfwwKQC223N6RpXN+/eyT6ZTdOUm2ZvF5C9cgcbFXDMKR
rGK1VkuTH+j7nuxVgNpe9k4qJnl0aqN5a300FxcJ5CleulMUzyiIbVidNIo6HfDz
BpsFi7iinRENex8FOtqQDhgEbEW3uSYbCHuu988flPGefnFJ1B76pYbMjVxmESTz
MJOQe/H+kb8njCugWcVsu98niExZSSKd0Dfv6j2/KxRmX2jZUAr3jjA5YKux4Ucz
DBsa3eaxpZ4brcuFJCJOMwSAgQfSGiN7Mm+OdF0gyRH3Fo2liX0bkbYvyyJA24cx
UvExoBAC0A1+lH93KmvkxKAgblY15E+venbq/Cs4W4FQbmm2zYC8/GJyeCZ+IWAq
89aS8RInEKsS30Zbl0CqpauAg7exsh0UivFyqL26KmDP/3n8roI64AtdPQSAP5qn
u0liW5iSiSy5S6VXzyXalcqTDH26ehXoIa/23i0h4FUvEQvU+Ws7YFamN2YFK20C
hY3FkjVaX7ELZ0TpNwhxsMlkwL6RuVkpjyvvl7+9cAXf+nUXp26mT4ipOYKSfhX/
bIj/He5jaGypMUa1hHuYsQp5LRQRvYzuZPcoj4PcSidSWhixF+19VmFqYUFkyZlO
TVa+v0XsRgOJPOu7dM7QweuPaHscWKjEsGQOWzsZ6Kmhqj5HYDpsyCJQT7tZx3MG
l70XHuKU4E0PgBzbj/DSaQfUHU+58qsRj01JR7B+Q1JI21IS41bGGWJnf+u5UqXk
xtqCDz3Xlyb0ptdK9I+czu3QJbyPsJr7s5mCGYZ92BajHEE+7QlHVIBRGWDqd3Cu
++/OJlZ1eJNzEnPGzdsVfuZzam5Xn1YAExMJYfiAbG2GUnBkR9P7oOwJI5rjaRs/
6wvewSfWiMTSjg8yZfGVV59HqdcCrGOm3xecZxQzD86f/jtGji1U4Hc5dbbjjdsL
tVH2ncFANVewKcIOK7apZmInq7KIty0XkXN2g7Ww4Zx5yiVPOS35aGopAS+did50
gmFi4oz3hsEPwLZTukGnpJBiCbXLjWn4acIXfJqXEWVjgkYnu1gwUhU2OkAeZ+w7
IYR6rCCvI1rUGSXkL4q8520B8c17Nd91u5tuhsfnjV7AdUsbLGJWux5YiYco3fB9
VERA1Z5BEaULxkgtj9S81K6xzqJsrbkLlrYTuTX6efq2tTXbVTz04wBAwwKGhPPW
vmt42gaE66mnj3U2qcxv7+3Uk4TcqgZ/E8Ckvayv3Es+ir7CNKNXBkbc1pTWUZSx
q8qqO4PqV4Wxf5Lf/yabeqphNQAaFqzdZiDVERS9NGibS5tYoBMpReYppviLLgNR
mqvSSre3ICfqHGpQaOe2+0mzO4IGaN7MgkJqoA0QAy1iz32Q5/4vv1SSjoLB0PGj
AOId6TJwBV3A/wfqWpddSKfv4NN9YeQuGH0etdwGHRCWjlPktcYSNw7QrY1ZwDLJ
8pf4um7AFPSX/USZ6me9ZTbsfatAGXGS/oSzKTiLz2VB4EPcVkL5aL1MuxzXjBcx
9aW+VBh/3HYeHbWruT2uDWSv1v1Crm5GxHCB5B/tZ7HnqC4tOTia8c6SNfsA1V3h
sR+qqvHa6YU1AMFj2WvClRnR7GI01T2cLzD52pve0dAmRwhxozoxHH+HHqh4uXzA
2+To6+s6IO/ajyEqnNSTUuAyyUJGBdHFYWARTPE5koeoC6aidSzVTp/WHHNQ9/1h
m1Gk5JaHIAsnBdMQ2eCjtewcGKtQaZeoqzlm7xW/u1CP5Bz1ezzs8pldSJFHumyv
TXS8tNd+A7/gffq4qFH6o6XWHsUm2pWBwRMBgrSGwCX0z3hFjAS2+vz+LhQSibhG
qQM0yadWGxcTuLPhs36iqEUtZuLvhG/ubjr2S1qTJsBwbEfWjtXX7D3ge9yF9ROn
Y51a6bwpjLwAUmO21J/xIISk3Okl3A+ufeJikLDMWkkZf7LHeKAVAM683geIavs3
I90koInCbfRB9ukBVLSvwuGCemDr0BTrGNApAbZTA+jlVjRBo/LZxbqzEnInHaeQ
3FSjROzP7sOgFCXnzqeDXd3XWRDyUbRdasVx/dfyp50scJ/3wvA8bLYy1gMRCGxM
HvG2o1itrs3jQcIiUUyAHE3PvTL7et7pa+jkCTXjl61318fAWqrHMOHs2wXbwesW
LPQpBMCDO/qU0QL/tnSkz2Rdvs5e9phRl1yAXNsc+E8KGFthAvhBlcMsR+pau0Xh
JA4VgXPYGN2CQ+M58TTFvd4o5hdwEfvlqNrvwahk9yjClqDbtgMJjMhBIrZwBtRD
VgyxAxL+YI5jD9xNImK9pYW6DENzMxSpWYPO1/ieakY8z/ATs49H8lnqS2xl+Rin
7VK7yukjGo3d8zk1DYPwv7hEEmqx7btMQFiARcrzPLSn191sowEIK8stRBi9NWmH
JMiR546dqD6dd4+6M1tZ1GihbLCgWQ91eXbfWRUbVGTt/Nbgk++9QQAwG60dGbQz
yLZKzU/1JDqipQLPPyzoyf2K3s8Hif5fCm1lZ0zpdBSoUVfy1e6EP8J/jMRNPgc7
WSb4s3tSe3kjW/nXWIcXHxGiO1UK9inrBAVEyNCqcK9OxknUNPj5vHFy5AA93VEE
OmZTUnW9aypuIVaPJW8tnneLd6Br435P+089cVx1R2nrLrVGIyCPX3uGS07R+mhQ
Jdd2W7mbnru1dt33W7swN4cdUVaUbjruqnom4b6eFhC8VRd2ySg9Zwy6pKNhuxE2
jw350SGgOIwfepzrRyAE+U04DGZfVWBA/7FpaeHiSbB20DxZA0fGhu/Dpb5sfGHo
U78wdY3br9r/i/pqI8I6HQt3W6Aeo272HFwqc63ot+wHyQoOuDaxf2WfTzjK9xzC
vuYtmyMzzGNm3D33SkCzepl50eqV/J2P3AggMijnjLX0LIrvjNy0y0rlMjMjoA9h
9Z1ictknA9NuYjFcVD5Hz4CRyrr3yEsTiPQm40ROAMRJEKWGxEmvsSP+CNKTvA7p
4Mv+sy7fbdMy5OuTE7tV2lwb9yoHBAMsCN/F8/QtC45a/qnGN6laMTbD5TB5HoSw
vZW4b7kpPwrICkagytN/eQ9HZA6u/fLkffLV8MmbXawBSMABkNSOUjVg/bwL6wju
i3DywtdadMwM8eZTKEswt9wnxf5/1KaC9XjnBHYdwgbZSNWyxn/7qfZ12KB4IUjW
eHHSDQ8zCiH+qsc4TyBcru7bR0K5Qad1QHP+3sduiS4oB2vpPqWDb11HMHrltY9U
+7RKW97GRiU4rF03tfSTX8vZlpNV+qJ7Sgb1S5JoXR+aEhEvQHS158KmWDttBC3w
5Ni0QaR2KQ24zxWBeqmAipBLAYabOictpOeQqTaPQr5TruNdAoYDdxLumRvyKfSw
e9XV9OCqWD4bDdkVFIPjlisPFF1c8ZGHVqG5qMUTOXoB8XC9zn+6cyZ9/DgUqliZ
5dXGNTAtLmI7o8SIyBVKsWaxG1gzCoLmTCgzLZkzLs6gZ5jrP7U7dP55Y/LhPgdn
3/QSBYZx0NzDfCMZnJrsg5ednmGtw+pxvUAHmZXnGr8zi1OymBkAemKxbLyoiyRc
i75kucUia5Qmk2Gm28+bNfl0vpc+WQ35Um58NEZYvx3sim1iG4lrGblpfi8v4071
AODYAe7+PvmBzpZB6Sfxp93eu+IZxKbAyITsvieDXtSyWeRKgqhzaepRXZN+HZdV
RPybcjkskHBwVr79C3HQMfqiw84GQJS6iDpnys+S3Hga8NUlJtXQBClmTcxFJ8NO
B0rLkFm5Wh+zN/zejvtnW+YsCcu8usvz/EzgUPwkbz+sa/Qu3fk5VYBUZBwv1Q7G
YeakhedNwmh7zhWB6Wq7IiDER/1sbrvS5UAxIfF0/wkuxiC2jiy7asSxItSU8Qj3
MBRFnPpRSp5ENAEYBEkkRcDf6Gher8ImSh1eGwlNwMUCLLtut+0+l0u4Rs3+61Sa
F6TVoSBfeRLHNydyVgLZQtfS3vT3Pq5V1G0YXEnTnA1dKrTj2+s8JASpMj/2MG0g
OwYbcmR8dwQUesDbHPB0+7hoIDa5dI5q8EGSA8VzMLTEis8lpnWajnJctZgO9nXJ
hxpoVC5lQCd+zwfgWRm79uTcoPZ4ei3RI4GRk0GmvStgS8sX5h1lqAxdPJzzlluo
6/Z+lgIxgzOfL5engHqcjgP6i8/BpXJDBw2mxH9SfUm1kL74K4W191fMM3jPbnij
3UW6nsuJ0zfUvuQv5gK2i7pcAeT0IcQ3FBz+YyCl5KiPriNTHRCteYZegnQlqWRT
6ul3eh2qO6fxU1/gVR1rqkBXKfhZnm4IwHb7lgqoa7REdrwqY/NxbVykGsDsrb5w
VFum2GWtr8ChbhYkV4v6Gy+XYqeHuSxrVRmnRkcBFwAUkCxugZqUX9YwuPn25d76
tF25/JJ0mjfqBwilWIWIEjr3l8IdFFtsQ3dON7lsEe0+99Izw/u2i173BLYsEkrg
EZKzkApgGox43lMtJP1Kdsx+nayjeo70bycHsFNmeAUecAKfbR6jtv6YXWNpOdeh
qpd4usLsdGuIzsEvBZ7FuxK8tIV1XkkR25C86+H5jJbcvuykOKRU5n7kXlsT5yWJ
dYC9Ao7JtsLgUHX23C6zgocf99wLwskBgP3wjwM2obNPzywKgfvmx4Br6hNOez7i
eeUDKmSLLAXXDJ/Jx9AyO0v+9oG+NLlzHiT23XO2699ddwNJOA2DqUyOrr59lVIh
RGpngQaax8QKp+hcKZzo0WxhKmX09bG7wUA2PMn/R9WTh2evT5weBlZyyTvVv+CV
H/7KlPggpspQ4fcHJtWSvIcYbN8adggrIYqPPSx+n+0wL7EfnO9BBOBK3nOzbObQ
7CdCn78FXmeMxTJcxZd5n/U/cJ9BCULQjsLArlz3GbJx/CUw2AHYSoex1qcHnmBC
ZtYB1zmkNKw5AFNtB04WP7vfVVxZeITp5kBg5uQ8JjsfqkE+85H4OWuw03AFQGY2
o7GPZDxt0H9r0d2Wec27FzXwzL/8pfbRCcmeYlLldHHWni+24+ds4wniX/FblGjf
zOszR1iFoBiB3OaIjsq5Cx11LJlZEhqd3UqszUUgn2kDASJzQxc/0AXG/oJc8E3R
YuXOj6KQ8cgRsjxIxSOvJvjxmzILfmnNpSUF9GeKvum5EI73Sm/mrTye5sqYhJPv
kglzX/mldA1IWSs6AmixGfECxotjOmQsd2EGQbZFFRQsOV2D+shQeqxE2siEET8S
Rp8Vw+hdplNnTlPP/DmzhOpRXTlxKUI56pSJ1MA3umAbgC8LMiC4NFWAPOdcpq4F
mv4FyWHcaRk8qBknr16JQogCq0iLQ1eOKCQ7SH4dFGCtk/YdgDb4Kqn9Xbc89R9p
62GCb8P+XE0VZfaW4mvYeIZsAqsJXGHp5E8Lbe3ljrl5h6HL4PJii83haMz7Tmwb
oJY9bWmx41zIw0vAYF+EFXePYH7EZIgIwGUABh1w/f99oolEdDcmGd1sRfpubHNr
KLZlaRnD0AqCqIqMCAWA0s57niNbmOyh4/MfbeKThwlYo80Mk7hgmhUuSLHombf3
fopGmyEN3ddC9eSwRyu1PuhbdsPbR5fIREzIW+SQ4XbHmTXb3uKVTjUV30Affmok
jIKtQQevJ/rSo+WVgIE5upVuO7vn/xDGhT2QEjARe506V2Q9oriE7ATYgnuLTtKq
dk0tF+h1bmFiA9qqm0d6otalRXsQE/UyTLEPuMbbS/SEkaeSyx3lmxf8mWFmbgex
k56RUobIy19GeEPFLr80LQ6A+rwHzUHP5y1UN7vNt8V5C1nhMGnxia6nhrSSkehl
jdzxg9ZxbBECYlKR6bIhOdl6gP9sDBH3bKS3AXrNf/uo3cDDdiisg/2EiB+3g884
1/FR6k9R2VkHhAFs1yZL6v4rQwnz/y3Cy3maOo1t6HWYM1ji84DzDTTD7cMRRTpY
0LonjtvdFKiCg2UzWAvEe+ACoTZ2qY1Y/rwfbG9hOX6wSglXQaHr/j7Fm54cVWAB
RMs9S1oI9ymOu9z3+HalbM25XPv7uetGTyVxRXh/q8yupZfK3wQFyO+K+az09pIn
4MyhKiQk7aag62qV33HOhzK36MlY5Im9X2qyhDlNBLOkuNnVe8wJQHtRN9fjmii1
4I9CUidGvcils4TqeUHBfmHpLhjosWpMgUwAwNmVH+YbmbsfeCTd4oU6jjK5vG5N
KqYblZYQRpj70a/DU6ZE5REBxXUZRE1EC35tuCJDSFbfafzttsXxtUMgHPUJM3Rx
6KOGlm3tNC7MVoKsnhsszn9PtUuMVRqBjWARKjNEkqzlINrQgM+J9jaA7U6KRgyL
6mzA/UvJiqlUIZxfzYSZ7gdCzFCFIa9/8IBYQ/Arcbtvq5juD/Cqpn4Ic5ttWn4P
naj4kTzxgy5Sy6R7bgmSsrdrLDhgJV9G9/s1Qb/oDGohIDOyhWVxBvUPblFghsGy
t0qYDbpQV8uSdxdFSQzQ5DtnbuOIOzdtjINUSWriTGr8a6EikTaBDwnUgKI5n0F9
UFILEwEFDoKu17DoMSXn8XJEHs1uSA5O1cG4EyJrOHeMOjnJjx4x5CPNTrfMuH/r
NkJXhlWqYnOKKTxqBTMcYMfwP1dqxUT97VpvoLLZ8n8iEPukuRKgghi+eZl7xVX4
pILkAQo3wPmt0ZEB5Lr/ix22FLmiOwDGzta1d3EYN4KKAuLakbPC/1BDFmcndIs8
hrlarMnUHSWiQzZVDnUqh8ljFBAIt1QbipCT9vjbvCSDkKYsqLjv1Kk/ib47zSCV
wSyo4FOVkXSjU9Exw9JsAubIeMArUf1lF7B+D6y2TzShcKn58xLJbfkfuw3KJ/hK
W3s7A240dDqO7BWD1DRNok1FGtPf9drw4ckZbYPWTVmRO95mKYwL4Y4RCd0RgECj
Nfu4+SbzqoCzeRFw62u97mmU9b6fpTFs2RhZt/tKSL9Bx2KE7RzZnfhdYSwpr8Mc
alUwjNpfGno5z+RGYJLQwbnk9B8cPARMjfNPHKWmqAxcnSDn8CyFtLGyZY5XdUZr
2moooyRtsyRWrPoEVW3qdxLpBgI6nZu+hiQ/7I++IIXr+PBAc3mBuoXW5d6N8JE1
Pp+iC3Ort9zCuhtaa9Iw0GslrC0oUxpxcmVywYaQ+kBYGpnriW9Li7jQ/+kvPdeB
ZisLw+0KclgJ7Y1VJltp+B2HbW8tPzZus7wJGOSnHgluHgUhcENk9LlgUlkWPmcT
lvcr+OfWBjX1AmUIASdLzuR9NvGxUCCLMTLCCFnUEX81hVwTvw7jhRjiNoTPrker
SxKzocLyvre07KxQAgnU24sY0cFyr7Z37momXtUjYaAibREZZxaoju1VgqyQtV5m
583qoh541A1hyfvPkfrgVUrEDB3Mmk1mHMIlAyHL5QRU7qOqYjmAxi+95MGibrNh
XhqXJD9oC8N+1939Ugr3f8jipZsjTAfLnHLUf1vQcqMGObGTNbyNgNZ7gzc8OgTU
Nixw3Yuu/MoWvS+OYtK9yJsMiyaTpOb7IGB0eN/CBpDAq/fHI3f42kO4DUSwj0Y5
XzNrsTRde0NhB1nNJngBrI2ImqntROi3kcr5EB3IkvhRdAyZihDjkiR9HVgCJQjg
EKiWFX/mPRduc6H+LW2MUemUBsCXKYc9BS532D7VWZjMMrqmCF5PNjpKRD8PCIOc
w8WQe45fsPEVR2OcoQRv9xTLs18Y0xHFQ7OapjD/IzkLBmVK9/4BQffEl9WkiaO2
IrAa3pCiiZLLwai8toDZTOxk2jmPyv9yZ0ReZpCzQUm+Y7B2BJZZ/BcbIsIkYzIr
jiIGepvoFdAP1l33rQXyG15jZvv++pdnz9EL3NiUBiF5by2StEe1FTR+neYOnRzg
clRoup7XiopVECYKifL3szew5g5vjGV2R0ryJIao20J0rr8Fb364RprkBsRW5hcY
rhJ9UNNyB/JomwCpIbPMsAe9U6uYmlRMi/xYVxSKeWFZVJWZKGz9PFYEuS80TYNq
CZUE6z+QlRLqJNuLl+C9Kacdyv//Zc/bpWWvyaiJazRu0y7Z6YPPhkGjr4dhuKwV
TXvt/2t1uAToUAN35NBtfitlYji2DDn3eHePjXN2BpDPlnLCLE/VWHHCZWCwSqNE
v3d9Pl4dY8Hg/14w8SdlN8Zvhj1IGnWRz/cda1SKdsTch6CY8lxvpgf8OGksWsla
gvxjTKX2+jKJOd0Cuq9mo2I17EY+vLWpyqrtky8uqVdgpfuv/CBf+NlLHOhpwmAE
3rOUJWZiFh3AItLrc21stbAARzxXtg7dyxMaLcntrF3/Az5BoOCKlmLYkoGtGCrx
fU8qrXo91rEGlbVrSgm2sEspF2onHLMYwqFQB1FvVQQ/AxKQtqy0YuKBB669PHh9
PXt+gyp6161p5IhwgPsUFvvPlqqJWPgt+ecsUPgcUCsBJHASVmbuxv6vFrlru7Gz
OcF0bv3zkCvWl0Ccqlw3J7JE/6ZF20yqH/khIPlEwTELZrMyJsx8faDmrsOKPmRy
vR4wK/5Zz1WTxV6cfYuszPNpQA3PfPxIKhJ47xF7/bJuS4YOZTW2c+NtaxdF7Gft
fBgP9RUAYVWePgnacYRxpYDXEgxBbLketjwFcOTTzBACakob8cIWH2gvjo/xwlxN
hhJ98Y2TzwmQ1Jd3LifOc46t2Z7bZ2rNlrj7N/f3M76XGJyG/4GR0Wn075fJRCrW
8dfG+1aH+/LS8Gd+J+CCDhFUAef4yU84oGDuhXIX4UxGRikmgkRzhyChumPeECGz
ZNc89CqtoNjM/qIhXne08iVDlun45beORy6xJJ7/bH6Y5ueoYwFAa3y4RsDIVnfk
rjuKL7kEt6mc+oWso03+P+d6eqfMxVrczAK1puedLmsERMaAkLMdZP7lD6KwfW0U
5t8MWsjHmYnozndNHEDxdQUBpsGTfOBv6CpA8FczXgJ843K3E7Gyj91Slz3xuX4A
nakIIsWdgN2plkq2sZbuDVSH8pLOyUZvIw9v0CdSFsX2c33CprMNR50l23tv4gt0
S4U86OngxXhhcBf6SISTaVa0XR3OUSLjXgBjiIvTUm5+jzdCgOKe+jij6OOzp/Sb
ONI8O9eD4lx806aFZO8STKdV1woXYHb3MSLtD+kfTQJDSxeSeY/E1K30xWrSaOq7
9DbsoKhSzkEktVMPb06L+0uqWtAtibdmCm/4zbGOLCL4F5ROqmrwMbofzl5VORNO
xu38vy6VaTakjcgNNf1aW3s6fXgj+jgFglYCRy+jt+Zn9tjjQfEjbm8Lie9eGTAo
1Cy/QhXX8r9V/75XdQKAXENExoM6y4DCOQO6rLjujAG4wq24Hvnfzn0/4GOi0N8N
2P5QdzWvxaj7XLFRw0izg+UpDkW39yKc1TjnEFJJhJOEJM7paS6fwETfs0Oeznwz
kQNh7d2SosLbea9lXYOJmGWh6DB4dSgCTO/VxW0BLDgQbFvtcac9QXC/S9XN2zcc
UD645e65edSeiOvTCoY5hIbtUz+EwrHMjUPOmrPuhZn+LA09NHOmssddX4ae23Cj
vVzxx7KwSP1UF6pYVfAZ0nN8BBScwg/PuwRnEyf1hqF0zYASsZdIDEYpWWE6cRD7
TOr9zP5UBcnBQlHndRTZvx0PPnemvlu8p3us2EeZLpV3ZeiX7yO14ZZln9I5IhtP
f68BM14ii3QGelMyVggeE9uMcTFGxvkS/e6uSZHtOLK4iSyh1y+5L5WbcyvQBBkj
JAO4C+dAnLsOSNkbG0S0yGdN7EzddZVt5FUXu0DLh6uLA/dCrzuY36L3tlm8ajke
L45J8JZIFOxMqLm+BeJjzhPkCrLeV9otMD8PG4mrSlDai5f5YAOvuSMVVRG6acPG
VuSpv9fDlBNVPs7vR8dqVjjRT3wttrVyc4uvLWStMV5kOPMoYOjYugV8IlZg3tlG
SdZc+MJPbgZb/fMmbpbYWnQFkjxg9YcoKGU/FWhgKE2IVw+hJnVYTaUYgEBRUVu0
NMLHlmFlxvwH8geYO5l4/IQ1JFemzfIypu4Vfv4PT/E9CzArfBC1nVrE4F1D2jMn
/7q5nUtOpiWLduzxJpw6vGI9GRoCoL18P150JnYyjYAtdDI0ZbPzeiuOGj/AmZep
HH0gAQr+GuQk/xA4G5NQqle6kgiQZ3liEZNOz8clgrRWQVWRI/tk2cboqh3ZwaTK
sk+5ld7ZpkTK4swzTpON0AU75oC64iV7ggnNz2ZqXLihSryOcc8/LYfZ4kK3qsf1
aZz5VFMGOtF+YDMuSF6zWVwnZfvcwZvLPQeZ2g+1NX+BgIoOAxTL0eUf2F1bzix1
YvJKgI1lpEWZEBLJK7WckrUVhNvs0Bti9eXBqzPWZY2FwfyoSnG9j9R3bY3mD3ax
6OovWgqzW5oB5uRQ1idB5Xm6jXbt0yOiNdRm+FYAiHGfukaifq9WF9Ak2H8napIu
s0YbUrKUDby6fKmSVq84BJWU1XARxXODGhyWJG9yUipkA7RegVy1L6yHBLeJKdlO
nExALXMAqTEuCMFx7j5wqnxGwT0ycAfDfQ7msM5NF/AVtGSfYLg8SdUFiZRZk+md
EgebotCOG6zsZeibHVMcaud/essczkfmBeWtUgpTA75xwdMv+gh7dEdmsbjzRylj
MY/yWYXkg2X4YHWH5B5087TD37tj1huAJOnMdrVU4qK+Syjeu78fHBgHxKHPxQTM
5T1UzuNcfkItveQmMmgcaDpl1JQ6aK+nBMpX0g4As5dr1o7Hlt85IPuNBSiDc/Gj
bNuUp3wbRqjXTLCTef3a149pS44/oqxOfhDMH6UyzQOBm6Vvf4EPi2+KzCuMYj7L
bpNuUL4Z1lZhrGv6lccWNDANq7HOOkWhcJ/Vwy9cQxyLdCNoLgzTX6EweANC993L
CMb/2ymfBNyZCDQx43Mq/vPCCYkYo4I78bQEVkyvViJvULMu3KDYc1tHYMiPbKeS
cWjO0ljoSmV0WhEblOYweQhk0mKJAfBzqawhDdALLCL+Ni2ZzDzCAFmDc5kTLTyv
Qix+Q/dqu3XK8X7xJHgCHfyoDVKudCoyFbwQxwnGbDKVs+RXk4bYGn71l7s+bM9w
LdnNe5VTwtafgCA+/ia4fhLgLp4IH9sVM2TquDBRAy9ImtS1dc+vy7jIfKMH/ybT
7ryUNgA1ePekLQv+8A9PnaDI5DmHHZ992QBKqOgB21ohrteI+jmiZVH1gaYLgJiI
rZ7zKm5yPYjmg8/TApR7qX+UMnn2CVzJ8bmYDBF5v25hEIv+BIk4S+N2GUIStirn
skY5D1kFsvXSuDfDvEMo8tSLMInznWU2NM0yBmNUGXxzixKx0aQgGS44ySgETOIm
AzAt2Q/SlyG8pQhtQqPouYa7TXcxpS0JjuAYMYWntzOzAZ34OB9KOC5Zfj4iZwM+
QO8XgqPgVu8IoeSDSQyggu++qa5pC4HkbfQrFVyJANGTVttSraAC2LQktBX7uxMC
Yb8EMYzOVkjmivB4vz4pZLK0R/A06DPbQYDtf1s0hos2UIwqQ7bDGbgVNn66DHqK
E6n0QuykK+zgHkYwWS9IElWUcp4NAVeBKKJ6syLlmRBZQmWH1ADbkUfZqQQh/Gwg
CbYeQ6aHtdkQKvvMq7TMMFb2WX7fjB/GRU+GVK6Zjl5DYdryWNzcDY4AzZznojAD
04BlnLZf8AUMreCF5c9xlr3A/SKRRkBUUAhId5R1JU7GBuFs1IzlR9bFX1LXP4Af
2MRcfcCRoiHHRYOCk72RxjmQI01KPWZ1iHmRs39THVUa1Ew0jh2hzW4Zh4+sTbog
lc+e2eDzCtyTdD0LgVomPtFOYJJZ+QIBBF/JMvwpgfClEztjCTv49Zo2wW9v0y27
i5sHGeqrkGoeeiVnDvIdbJ0mNoeoMNtdP1K++tdHbgiT0F6ugMYRo/NGSFEe6jAk
x0y7+yji5l7L3bYEPGz0UaoLc/j36erQDUypKdb3xnP/RAmmJfwqSgI+VX/Zz/z/
Np2VxyC47mQVQetIWyCtIDCYMKPwaZ75lZ2JAbWWrkUaRCd+hCTcDqppw8lF2xfA
qW5wyuteyxvh2xn57diopHDfKfFaANx2CAYRwkSdVBFdRJk5HQcik9mFKC/uqzvd
vSGUNsiQFdiWyUglqfs59aHRyjUg0SUvp29TBUs62LBDrB6vFYQ7mSn5UkBPN0qf
KoHo2D3IcRrvnGeIWy9TCaTCerzlZARH/7+g0sRjB0ja6cky9k9xf7CqrlrfZ/wi
1fyRV7YCMDF+TgSv2xrhKmSlRb7sGmF8oIepMJuWdIeZjaLtQJn9P3id12ng/RT1
AG/eff5aLEQ+eImPvCR6eG/9dRI4r1dmrKPWksW4BfujDMzcYedRXwPyIxJU6xgj
RJBExbWTEyRbRya9JQHkcbrHvmxDLoDIgSJeJvfdf+VyvQ659DMCR3ZMKKqQzX+o
bTLPvk59WZRQIJ681lgNJqxjbQHan9WUfuTVuO7LK8usSIf+Kv6UOxniC/IJjd67
zwuXftU4GNl3EXsDRwUKwWYYYzgAvOfxAQY0pfkrqPyE2SkOYK2FuxxS4XDj0IzX
0nnq5E/ztUHnWahICFKROVxazflnZPtYw01BwT2d2j0L9UV5rFJqrqFYMUG84Rot
YOV+g6D+9zfzOKwhuUoOw73bjqZCVtYqRgqP8JbQmgGTU9PsxvcrXH1nRL7cyGrN
cFAkSiXy+yMCew+S5d1ik3hAW+IJDT6XlaVqsfkIFUXlFHGATizYFEWc+7iyejxr
qXKq2o9i2vU3j9Op1jUPrNnkinW16u3ekR+5VgPpt9EOvLCSyGcy9Tq9e/5aszg4
ibuZG/Du45Y8AsJUC6useMUswXVYf7yej9z91SjeE7rbSe0rIDJBwT2ce1tT2k5x
ht4heK1Ktg+AGwdiK+36OGNixq6fBpbrlA/zGODeMFlz1WoDlJkZXokbIUACpYkd
woh6OzUrAt29jLXrRtwivPWKJj20E6BZgbhi7oltxl13wCzlje5thxhS3KK6TnmA
s/DsMaFiGwy9VhHmCTZy6CjCF6uFcbWtpoShcwh25uPbzWi1I/y6QsmU+3//nqN4
1zm7FZkaanCdJQvQ/w+lAOkyszIg2aFPR46zZo6DbjwZRfOkn3svRJ8GqQii22Yd
xNH0nRi7mjdmPljqG45dCG3XreUV3yLN4yjxg6WUGYSRYOaqROy8uX6HoxNh6cPj
DpB1RLnEQZcHduMRCnEyqaGdonfpgbPF3HFcqtrqIuq+rZoKYJH6XJu9yUa0xLtz
MQAb3iItSXFuPzWzVAhcmRT18zFPodBl+SiiELy/ON9kiSfZRafWhko0vl8weoTg
IXYk9QcWcwKEfB4Efj7MGqoniWauIdux580gtJVjsOlK3Dtj8M8znPKXv0fh7Yia
hDEpfWdVFE8J5eCm3i8KhQygywFnR3oNZ0y9+/zsIb9QALUTc1FqWTSSgrpA9t8N
o2vojBn4jsM6LTgqjGdR1/u8xUUElK2UuGnSU7TEJr+lxhid2DGbWYcDV9l0mKPV
U8myW/fb94QMNxUwwzL6w6bYrsOzl/bg9gYFlYDvOjUwpoOURd0St5CydHAmqeYF
XKuCwgWwPNnFZO1wZjGU2fpJH+CnkuVNB8sDzK3CMyraulfV3Swi42BaVJ/d1b6S
Fexo4tRlG2Xy/7CMWcBao4QBMfHXkttKLEGIxnvq7CxnfrN220cz2qwfrIP806Z3
41wA2VvXkDTQwZtS10wFI8fVPK6Hpv+bU7OdI5/uBC8y9b01AdM+S7csI2mtE3Hk
F63A4aTLQZNWnwFPvLwdBnRg0inO4ESFmFQsPxiwizL0jcqrBTYE3eO4OzyXFDJD
TgItQUGCpV95/2LFcFZPllgAX4RyWj561GqIlWvuiCtI8mcEwIROxR4P7W302jtm
3/MvFZ0kACdCfu6HhxIPl9n4PROzumd92PQrcTb9YRD3hZaA1+AmVC1vCUT37DBS
Dhaz0H2uNGuYADPg+H6hlCxDxgx+7fD7OljGHWT4P2Clq3XLG+jg9MOtErWBXvEI
RlHnjFc0DYui76S+hJ7br1ajSOROAFePEfMt/Zki48JasC0JV2QQ6mSM0vP89HSN
zg+Qbeud6NEsQsREaYn0ZLFeaJB+El4AeSMP06lCIdvTZFUx8//SlTQ4t0+liW59
wmRzRNGTIH4BQCwf9eyHBzsRZGs6Xb2WWw1lrkFiboC4NfCNwPGinVM8eCvkANoY
i6Vewg47FVlZBm1zffQwHMHoR8MqnuQOUjJAEGdH7+aAJr6NVfgaA1z4pOuQDqzT
BSyiRn1qd0caaVcuXw1op1kqT/5U6b+5AJR9Jle0Yx7J/Vb/bp30eIhzaLt+NK8o
BgErPtI5iyK1qZsN4gAsmXXnLAGgn/0Rdkl1HP4/1ZoJ7x9n7Rb0r1mQh3ip9Z4O
JsTYpNDxlAoZHxmCBDuqjBICVgRl6DsDBet/zytkqJoYK7c08vjoXX0ni2oBUpU8
EUgOdYC9OPF5wIAi7a6uvPryh4jJC/ITmHTtclt2zLwhOx/UC6cxwEnZttkBG/LR
IIUSQyUPev4K60LQNVEjToSUPOQdRKClM+s8JkJzFP7+3cOoBoe1ZnOJ7Gjdi57A
iaLJVAiP5pKnWwBBKszbk759iRHDvB8GZuQ1uuEB6uyzpUSWkBJN1TqpTN5d2Rnb
9wIs9vC3FSPCLC1OqE8+H6J39x+ofPHbdxFMQMlETS0Yo+btcapV/tk536Bdp04Q
R3x21aFJRzemnS5GUNuu0JIp20ufrVqbvzIElwXAqnD0pK1d80kWT7m4KX5Zcy0j
LQ2/A4Kmeqn3Fr27D7X+ZZb/sIfSqJrHbYfjzh9SQah2BJSWkCcoa9eQsoo2Aa6h
PRnCCwLzvMmUgzqrENzpIq1GMLDYMiYOq4OS1cO6XE6vHNj+XwfvE5VPX5P/Iwb8
2H2fNbRiBgP1PpBu2F3sgC/jeh9vVySF6Dd4TPYfgHd70IYZ29lJbLb+7Rlam2YT
nIz5OG77Acbp4OPPwSKXGOWA6XKgCSYm8frm7oWUlB5WCnOzY9T+vcy93vLbT9z8
bR9LBN5Onkt8sB5c4WN4HB3SvhHHL8n/pvNzGgB9xTA8OQYERYBlWklVHCiCeq0a
Cu/ExIEGSk+s609+0dpFL+29HnyN+YM8CKCXEOxbB9o/fxxYwNyYS+L0ipsbjCqb
h1aNWDX8n+Ib4dHG2fK5hLl6rN4hKYSU8otUYZVACUtrEkfh9dsIS94RFwTlMyGK
zgeKibNXkMgjzeEpTw0plxpqyxcTvSKE5spoPYw9ppYV4DH4gjr6NHxlU3PVLTeC
/sOf87shhiSSlPRGtsJq82u+pxX8OaMmti1LHfEsaV4BFF2GLGsoLJSMYwaSSbj6
9uoGrqltdvPBh7cKY5e8FypBEFxPo0D+k6naxHu5TLD5RA1RsixaGupndWYSI2Hy
wJT1z3XD1pF+OBUjInxlBUhGeLXPjh4hOHeMZKTg6r6sGz8+spXFDj0wsbw5Oeiw
ilnYS8fGIa4h0mXFqi7J/HtUF6vN+r474HrNPjPDfyJh7lNEDotZMRsmdUZJu7q0
G/6bWHpyk88I6j6yZ7RdPTKMLz79kbJ8xLExu9EAr/nNX4v+w+asLe714SdZJQ1t
mRdlownKd9R9/z7cm7oPvk1IU5TYdsfRJJZZGy6R3zswzvCUBYbfECZVvg1TdJrU
EEWDPRWIZ8S3rFTYsm5dd/VDYGJCYJeuVzFrPm0Yi23y+HkMX1kCOiPxZ5Qd85w6
FneDaqoVFd4gQzgbR89ix6gtVLy5a2kEIgoXyjowflzSzXyp5pCIjCKuGl21PlO+
po2Lp4QX1TcMBw5XA+C3655WLlCaYYlOcQRPh3A6eWk/zomZm5ttdulIMu9ZxImi
g60oX65AcJw+tSMjDLqFCUc3uSp6bVJR6WVycpuOfjdkCgBwdnLt2JzwV7Mvqam9
46LqpZ7kxROR/vhCvG9fedE00WO4m2Q+qOvziJeYb1aJcVOjQ/iR+mC5LHwQLU4f
ZDUUF91ubsX/HFpvNnZ6N1QqMAAuzBeWj4cJVb2HGhtWeQphR0zGa7jPfxfrA0Rr
SgfwrTUMFkDxXBmAm5CQT1aUxPWfxkWL4/J6bzpIWMNwbWq6v852gtQmxor+KS0Y
2eHPmLDiEy+mZgLVkwhouP0fuQ7YQ8y+firvjYj6mSMnXUvGXjhM/ycwIkORRz3E
JIwKkzhcKilbnZ2ZLiLNqcSYbWGUlfoRr4tR8rcCkkq7qhiegfLjhbSOD+Juy9KP
FcYFzKvTxyUwUunmIovlPRB2B9TlkbPmB+HeMSM0z7Gg25OOFblWhJltp7zP/3F4
aMco5i7VY4FK41IgS9LUiyM9GWvU64eidV75LOzET0XdHQfZXCCkRSnyyCv4icvk
nz5fc2zU0rDBgvljZW63HTByDUjeaTH00uhh7tXkFMHIi9Y46kS8sLNd+1WwlZhY
PKOFJ6JsH6j7k0Kf7mLMHG0k3e5EnuGHJWGha5v5ovoqwGD4WW+sEUFu3f6kS6z7
cGC6sd5Sj/g0unwhqpFRbYZrBLq5wN2qNIvNCeY1Z+VDvopEb5gVlOLL7MxAetGn
DI+HyDJGlyFHAhH9izvDcQHBqHYiVZBM7NyWeTh+JUWhn7oZt9Ht62PjXkkoE/UM
gD5nP4RSdj+bsVGb0z6SH7Az57zxkcaMOtXXEX1GqQje1uIkAftH+8OdqcVdA6QH
PhWnBLFymk/x4nVnJSzXjgzd9DYaJv/qKbtfdMngZZsVbN6OVZNK4Gm2US8E4HOd
1ChYic4hGAJ36tc3DGZmxks0VwKI/KBriqcqE3au0lSrEeTooapGzvo2aXUqlDpR
h+t3rQuqn9zDk7J/mXJ8XbtDHhVzwotYiWAFxRJ6iku3187DJxMaY+DXCLdBM/eO
vyj0qu4ipPqiMnCgV3qDhv7ZREzKPcF6LWMSoGaNwHkkPFsXdV5GMzFw/rwarLd3
pYcMLjQImOPfmu9HWWudV15ChV/VQsdgEn3RB9mE4y7Eo8PQsG3VXtlDdUJfu1iY
QNuAeZ92V26xNWR/bNJAXiqPa5Ui3rOlsFfTlCTqHtrrQwJYhnlaB/2kyRo8O0lX
Z+6Am9kJgMGpAv6OOs5HCMt4pqa/2TSzzM71l1IbVONXiQ/HQyC+25gLes61tW1V
gCz7iLd9cRJJmz+OrF6+ncrcdLdH1CnInVyE0uRCYYu87vmThcpaXrf0yPfipZ0I
FCrzAOutZguF3A++ISfBFWR56eo6aeeaNpg8rpNb1dZPlc4W9zXc0sK4crSR4Zfa
VqQ+st5ZfS19DrPq9wn3Q3j+JigJW+i2cE3EZU94hf4RAnDGrH30VUfgRRO0xGhz
fNaxOJrTiGJHlcFEllnZ+1AFaWITlDMcRbvNVD4m7A+/qf2CLjpbgrf4HrJiGs+6
idp08dfQlOZm0ex+ZjhkaagSPs80y9s/KbZWMoSbJk9dSiP78l6jzGVD6D49dWGz
784VcrZwOPoDmh2/puBms1Qd1hhWsspCsNFwiCYas8luKYIP5NE00sSLBqbTEaLA
919f+y5eJIiTXulqDMSBuoABZZhKj8kSRoKvbtw0e2zsi1TJKw12JhxAkLxLvQq7
dqbimyFlaIg/niLYwdYi2hjDEXh8cg80cCDYDt9k+xLKITPGLq1oQGU3L/1zgdWA
tBXTgy5oHKSJYq5b60HjQwoShQHn8BBQAiWDdWU3P8BnDPz9UypLuhgawg5cKElC
gXA2mVzQB/dGtvoKOwFGQX3qfISVa8BJ9XXiiQwiiTsem9+BxxRY561aCjG1LGlR
d5v3N2xBjgpyol71cSvGo8fvdlIIQsWKV3G4JZ8cAnHK9KjIgwFh8Yt/GnE6rzbt
1ILo+PIq78EeM2Ki5WYq2RAHZzYJduwZTBJBCoqPDa0V9UPnnItyrV4kEo75WE0Z
he6MuyQ4ppAfn7NwNJK2CY3L2E5g8pknac92qqhpTKmsjJ1+7jZXQlr+fKsekVhY
1Ucj4grQ8gAF6GC9s0tJ1+8TyBgCafhRq8SVQDoz/S8RMmcI/BoZdPe8Qo80fj6z
T49S/I/k20NApdZUgolOw2HZptuYQ8xunWiZpV7a4BqniDu597/fwy6g0qhNGJQn
XJHH24YJ4BFqEIpTWV8NyT197FO/pEgPRCN0zbcmU+OfSypal7xhroINVAGjeFi9
XZLICO/QLoV3Ymd41y79mwqSf2r5omTLR0Caz6R4cggGYtV57h3GRvoBHMvUSICh
hMqUsCqiAr036ayV63SDQvDy+Uz/wYJplkCy+BJRr/e6VM6KCS9YfTV6QtSoXXNd
Q348XBf2qUZHKqQjSfl5ytZ9lWBdV1WxfuWtkvsKkbs9KgLWjKxLq3vfYX4sIpSI
DDcDv5ctoJ7lC+UEcB2ecPe0bGdOqHzdFxin4XPLLdshq6s9CSdOGlvLPeAXKP0p
lNS852IRMzLb3wEI8MuwQSlmVkgZjZSzpwCHVralkZ1FkRLbYgbb7OBxwmnu/L6x
Zh4v4Qzo1M+jYWhrqX2+HG8D42Hq2B8vCwgTG8rFWD200PaP/VURewG5fr73hmcx
jdjzyNBb7SucNRusVSO1kLq/xUi3Y0NPOu8t+gA7tDPzXNfIJYo3IMBMYZSQJ2NQ
bhl51kyTLUcwe/8ajf5urW8Ao5KSm9WifVYt5kOVuq7h1+4VwKuWL62L27XhHnDW
DmkNVS3Ow0IGEn1x6FzOii0AbjQNHSdYkFe1O6MbH1JySkh4HdQAMT0PVr/0nQmT
KNPGMNzpRvK1SPfctKVN4OnECNiggv0isTPsNEZ1HHUcJxs4PU0Msvby84xnp71X
J3tqx++GOkfkHp96SQnt7LuQGBnlAwKl0FIEedDqJ+HYRgyl80IPXtW/iPPZ1j7e
oFKqkYAWtjHoc+IM7VCL4vAdrc+6nbrjuYJ6/JA4KCi1EV6G/urdrIxhyN+EmRzZ
lVJ+LPITIAKQ3KoEKnEwlBe6YJNAoI0DcIATUWIHoj11dp4SLy64uPtEA8Hkj/vz
shYycyQPtl8yPVvGk+zSPuApmBtPfMngm85/5Bg7/Ua/EBErJoSSG5U+Rto1z6vd
95q1ikwqDnnSiR2mi55kilD4NcrpyUEge3vs/GPvrdv4kL52YeWfVCugFBiJmgmH
9pQBxr+gNyPU/EgN40Uq/i99A+/1XSFnR0sk2OSNE+XkR5R8qKPjIOqKmtfni1nw
UKcVR4mKgxhMQ1W/ab9YlHnNavHKa7lLC5jFIw2MxwSXq1lTkdMJQte+kYBJ9Dtf
B/z8ZgvG/Ouos08ladhg8pQvPKq+Y/8FwbMrHpZXVv6hPp7x5GzZUxJl5XOShsn4
7od6As2SFQJwQaz+LnhEvB5cOlfYaGJXohQarrldUo1c9V6exeiDf0UiOJRR8lGM
ROXB59gKfRQAKyBQJr49s37NoBIjBOmjqsulRQhhB+mKAhv4R3LuqMRm2AI3zrQY
rE6kP+CljjIPB2J5OkxIQEuu9waulKy3AnNakqAsbaF1/vZniABmaNvfO46T1oEd
cvMg6NRl0pyMZoejUIyV85dF+tn8ReBWcg4LmAFG1VN6mc+LrsF2sxGVGmCeix8O
7mTj/qzl28gx+FgKtRTFIWsfd8BtbpuiTVrz7fAqZD89j/6yUDCWt8pcUGQrKyij
mRa3cZeBrJATxaEOipEY1Omp1FQEcc0Cc1a3IjqT64qyqxm90uc4LQxoJUflu3kw
HSZwEby2aHxurA7uVXe6kU+FxhP6rbSbtmgHSllnQ8L4C92IcT8dEo/q1u3amK4r
vIfQP/fJV7eseqFbQwdKNeMBUp7XhBqZD+j6VZ9TfMND/ZEmwI2GjpvzF2b+svx6
JSt1KqXgEg+2vfSBFiuRRuiQQKSg6VWKH/zE/ETJ4oIgMqVQxRrWvRO85ojwPkz3
tnQpZ60KO+VJ/roSZJkLS/tI5HPeXmIUxVA4ihOuASM+w1AfyFA51PXN68vrBkHG
/KSaQJecOmyVYfCdXVErxDXiyjfSgqyx29An6SHbRId4evs6QXiiQxfFT7PpOd0j
7zmXpvD9gHP0yI7rXTc3c+/UwgFXCPT34DHfTFMybJ1plBDE2fG+UKNqzJksouXI
Zq5wElHKODPkO3hCtMRAo/CCXE3cZmJmtztZ59x9s4gF2CvUX/jNsX/arDnbBz0k
s2CBd83tBjWxj62VscZUo8QlD/LsK9P97dnVyG6d+Cyns1N0fMqGtC0wADpRkkNO
5/hDWd9L/Po7k+k4Cfq3ov7xDG6QmQjpClg3Jwe5EItg0Pqq6gpWk7u7bNJq/owU
x8yqxmozn/F0lao4fF2VY2HUwowCE7ctKfQeESODv06XekdW1MpvAfpWddDIP7Eh
ogDU0Skh48PEOiR2OwwOQPXNNOHEzeZtiWH1zkgMuHR0hXGtTzEP/ozN89MnifOw
+jNCYF3kSBSZhHkMhO+8ZBWqRJIEyb9m7b1nU2tIw4YvyfWCLDQ7xWuJ719GXkfu
fG3VBS9VmomvzlHvFvlif6JosPBO92EKNZ/u2f7W1+NkNM97ZQBPuWyt88/OnLuy
JK5PpVYW3Dbiw6PRtL74VPg/AH/H8Y7Nqx8QQpfIeu4W/hpfYY3uKlJYpRAvDRZx
Osh4SK03mRJjqJZGxRNi1LexK3y5/bSnwqKGAYH8el0ywbDYGTeAL655dXsY53aA
TOG1j71iYrEiQtzNk5LPjdYkWOIrB+dQ/fUXrJ69g+ddZKT1vkzZIZ0/9IQXtIOm
jIUPfDwxpMGqTZOREmuzclpF7oHGp6Euo8Pj+r7CRZXEjqceZYDacGVU2OlD3krr
PmEs9XlaC52rJZmMjAul17/W+Qq9+UVw8XKH/z5oxYJYY5m2BRZqf9E4RdwC738y
uT3HixhR/jyrJBPG2LN8fL5W/d4S9H6+YrXpTNL51A9SgAZwgvCPrbWwIAP82Pqb
UfHB9Bsqv8mrfJ7U9w1TVwPazFnq6p09fMBVpIrLqmb/JBUUhyBsqshtQK6vDy8K
198v+9HEn2wxP19Z66p3yMpIwUmOfUBtaqyaDi7/5005Ki2Nf7M9xzOBOvZFF4s2
akdshSTYaDgV2yvdp2WXD/3BDW1DjPtF1DuS/9y1N0YFSpUWUn7PMQeLRhlw3zpq
PjQRuIkf46daFwp1ckddwq93bHvcgu9LsdxXuxfEDXyhPD90Z0t7V7hDcmM4QEgK
du7vIlvUdZNx8evC/+rukg7cnuC/RyBxBfGvWI0JYcfRuseWE+7nTb+Uli3RFtNi
/7ZLcMN6/C/38juERoSKY3xsXl1m2OyOW/+c9rM/in4vqxs2oZGMcufdBrXZVaDM
zpymtV4Hy3Altwqf/uD1hHGmDCLWyNVVIXmLe1DHV08Y6igvCf2q6YR8HNJi+N1R
O/ZC4+NYU+RsDWSFKLW3yYptD1YbJLGyFK8xfkHTt5QcWAC90FdOfkiNb9tFcHyM
AO55ZlbAfIS1ElsLDWo1XwlDRl6Iu46a6lInPlF9DCkNwy6BJy4uQKdkYavofcqh
1Z7DdvUdOcDE1+8Cgkszqi77Mlep/472wQejWWe0vChDjVCRh3ZaSRZTQRKPOI+Z
vjN6yoCsEYUvodq3FDC3yeLIg4d/oiqBsQ/R1zsFdx4/iZDDlfxlZpJ1+JFfFqdH
a/clz0KXKCxCB2lZQ9a+3QBkqkUzCOW+7r8W0ROpKFalUM7eUobLSvdKdj/9yDqI
lMeGN/HJ66hseVq2gkPEd0MogFi0at/4+DX92ShVukM0kepOn7lkyCp/abYhCMLd
3D1d7Bx/nLfCVm2yMjhXO4H6yYAvI8+DTNGCpRZFkzjyGSBi0X+UXXhJNbSyPiZF
ltlzUvUteWtWn4GdlCTfP/8TCBp1D8yFuF4WKg+1S0i6DlQx6J0zWym4DYbWTFWm
wkwwSfGXeuzxriShH/UkoL1JCbagazm0XkH0dMcRbHdrU+Cu+Ajx7s4twXvOxZqd
lJyozOAdPlTG4HRikgUZPRZxqG3DTWf/dxkcKRsj+CSJ4RXX8GgpprhUYV5I75pn
HixEWe3cO+j2EZYuvX9fH7SPnGjF6OPLoAvGT1zNqOr6NU4DeJgqWS0qNCrGucCe
7aLsed9xEo73K74Ov+A7TMuK+Rw9BfS7gy7jhbBL4yRNeh1TuUmxafYuPnxZd7+U
LwEcdamP86KM5WBFMQk4uxczSOBJH1o2OdKn+VjctY/U1WkTswv4u3VPlXuZmek0
/3Oh/WekgNySSn960uSLoS2YolJFOtvRgk75OkRzrS4F9vd9nSbTUtjHInNpKgbw
C/UIBtoEZE/uIV0qHOBoUV3AAxLBk8z49kVULxZ5cw3RavLz3UFj0LUIXv2XaIHO
2qy7butzwql7QFAK4Fs6Wugqw+HPZ7Nqk/SKHjGYTV6afGVCN5k7oSY8sjKFy8TP
Xz+18BQLw+CAyWYUQNez2Ct9pKApEOHoq9XExtNaSZcrEO+xeupoAvr3h7ryqUdL
NSPHngWDPVhi/NwyR15Fw+plD+hmYLP77br8OyXEHMyllNpqQFKf4uFI6EjWEsF0
J/zJgQTBRNaxKjv+GO229J+e1ulR3npx5FYl3QngAP4dUclihYjn1hxbeQpA7Dtm
HFf4N6NKkhmVkXa5lgtYtakFK73ceYo88eHqGSZsnzAQZrM36+O3yKKz5z/USWyl
QYvV1oSMKT/f5McmPk2KA/TEEwdZaj8PEgAMwH8ccp8Za0UJq6DRB8YwV86mCWWK
6P3srtHaRLE2eEsKDh9VfVuGox6blJtdzhwZM2gBtIvf15tobCoV21N0RFfEn3rZ
6AF7lcm0oPLztUvWgamugf7DZOPUdhQFbD4hmkWBAb21zUlq0tujxzQt3zJp+1kB
6lNaV6mPLRIpkxxLUaVWX+pmW1U9OoxKUBisKEyoB8Erau7gRFQz68XlscYi/eSE
1ANFhMS0oivpuy0sQ3EkY1bTYZWIF8qKiN5P8Abw9jKEp2BhcS0QzVlGJ4UsX1tG
xHgFtb/erLMv4OaZiVB6tZq2bgnFrfn5mBzzZPzCZcmeEQf3tuRdefnHgzQKuGKp
ketAdfHmv3rkc4SXdTvU54aN05VfSQLpnyCsqNcZaGJzXohIqIe52/AX0sQCDl7m
S+FijSCSiBEyxIIPt9qMNfNBSf+qrvf12IpfK1yPObn8batA5TbZ9CUlEr3TzgXi
/FSMszP4xWsVbqtxYppJVO1o0zlduCu6ZKOGZZzfIRFX9GPydBMIT9punRk1IJDI
0h+cGHQvUMoOANayDyZO/4xTFcS10n/hIWGG0MnMPVqfA2PUDs8ugFJ2JKyhb3VN
Fcls5ohhx0kaYKS7+vdVOHGHYtms7pQ47jcWjhEgpB57ZsQt30JG9t/bIfQvOYf1
9bdBhd1WLprWtD9o0qswGDlGQM8avFmm1VQ9sXIkRkzYMlKY9Bki4Wa5zRjguebh
EnQ0135I+cOTaU5gbC6n1acCOHnDlFLKuLz2d2XAN+8QpF3iGEvSUaLZ+EMj4Hno
VPIDREjgS2vFVzZBVHxbt/IMiJ2efpwO3E4v1rO+NnW3TAPMDyvmvaMe+YjwAz+G
Oz8fbPJmcIHcMRSEUWgAyeesMWt4NiZK8dwO/9i87g1knQCbc0I+E3indSny74UX
ON+cgiB78Vpg/gsQ1pDwiPs5mLXSw86kp46J9OHhWw76by0IepXVfCTzPVl5wsGQ
FyIEYvyOlSD9VDjIDvbRVUixT9U4HN6Qkuiic/aQifLGYBfNRGrviFgrTCfMt/Uf
ELLoyfPoBEFcqKHnin7n+Qrccws3KhqpTVtyaTBvalkRBAs5sLi4j4jKrbX7GHZf
f6y7Utsb6AQqR8FhGEwki8fWlY+/b5dCyj3ApdOnPq5uzSf46NUyVvqtdczCt11t
PdgMXbGjoJ10Ne4e34mxh9Zpf4lj2OV75N8Q5iOUyfdTU+rlsmiuilgExl/yrQZ+
HaxI2jWqRaiSi5pAB9LWBU869oo3OBER7AipNmWRCO5IZWYEIBLSIdXhUFR7AkT6
QV87lVATVHzDSNvRqGaQK8N1YLGpH8GldPblrHS5vyl/3ZMP7PRqjbOA5JA5tZta
l0ki0L1BW1KrQazoQntBR7A//61D8hvz2t40nfqPrQQrv9/P5enrgXwqb9p1nt14
bEQuDrPCrj0QMqK/DEuD4d3ZGwK5q49VdTJbIARbKb9KcWf6xLh29n5uPI3ZWBBJ
GYIlnMAAzhcRqa4uCw++IGVdyrqBSyRl979SbFyhpflH6nv9+5zKI8p98ppCxnuR
Pk7DyLC7KWAeZuXgXAi7DTxJj7x04OJpEA3k3+K8fWYNG7/7Tl3LJQLhHWXiDCvX
6jTn8XTA2Gg6hAb5jH1rV1S/wVwUToB3CRcU+WanWkMTrtJUC6iJYAzgmfKOQgyv
BXFZVwfZa31VK2UOYyhejEHarZuWv05jtKhVw+6r5UHYFiNUuKK2Q6GlReXcpdu/
UVkqp61Odmq8DRCcKaHSIrX7GecaJlVCcKE9JfrhruUWx118gx5uIkBTiSpXYaoc
ZBfpJ2CAqR1QcFZ80rkunpFQdlHL20GP/0v3QKKACWgF+fCLpgqKkcnHTG6ouu+q
ltxAiNN31A3ItuRPdve/M6xwcae5AZ4a3OO4X3Qe2wS7OTCPO9yprsEL/Zpri4cz
lbvHZKPyWS7/DgbXdqxYQ6Vf40ylPoZyIYUPNNc18AJC96f/3TH93z7kF3c8f+i0
f2OXEHItmjETgTY2si6mbUnfTO6mtt7oLgqN78yhwWCtvNqnB2VzvMO8z/gTnT2A
yNpsO4LGwDT2/D4MAFk2CFxA+XBhm8wkRfYD2fg+YNFd4tjvUKuKABLmX2sJw6xs
FZjGkmqiBtrKLdZZXqYupWZy3sN0MOfXEVFpW511K0KgL+G1CMM2yk559Fy5Sovx
z0sZHR9XRZ2/Y+1QuX67L11nEkhRt+Ki6BuQiV4/dTR2KqKVmygFK3wjhBo7mTYE
TQKTkhGYxVTt1MF3gtCbYgGBOdA92YlA8WcQjxCJ3JPf4oMnWy2RUTy9wL0OsI4A
NZDJdeeh7jyM0sJ8DSmjceAite4MmgMY3nM2NNUJFJ+pvh9inbW4SUegnJ1W5A2F
XmHkqITkSFtC3tzl1fdB7Mq7izTRLeEJ16q/XQVj7u5FAzJS8Z6xzo2s8BveZkZU
DcVNjR1a92JSsIGwKX35pbkPKEXwKoeqXzd5oebuY+geYYMCTpzmns0j29XHoSic
3a0s8J4QEWli9Uk7IF21IM2Pisq84Yz3sNzOJdRCQDHSb41I7+3lVpgq8qv6J6yC
tUkDG0aGgN59/AnpG3th6CPreHIqcaO/8ScAZiSOUVX0Pnp7wP0HWAO4yNX3QgTK
Jj3nyaawLrtC3U/DPYcCaCzYSrgtUQlZUvH7+8psF+myyLYajzN8yy5EPceSDyPY
x5Lp7D57m8elZLXVK6szZI51yMPUde85pCc8eyUafASo7x3CRrdd/R8JOYM0R9ym
CHYVuWD6rk+vdFtl1PX13yOyyfql+236sZ/sPTCAQwRUlY+WJYIae8cN3QTl3JP8
p4b1JvMUloRKq9Btz9lin8fCxoQPiNt7SOSkHTb2S1pP8m6Erph7AzjSTbQHNgtD
tU6QCiRiIk1t+rVXQL7Hl1rPeXOZgxrXX4ekEgGNQxWUylnzV8/Q0fW3T7s8Di5F
zmwVCVrwbOgvF2vhPFOWTaZ8zTB8U0/mklrIqB4f4NKsKkv4qkUQrjEbDKD/TA19
QbMrx93tCbDiwkHuMSloB3d9B/LOflKQfR+6kM4iWyq6I2Wf+wa78JERVYM1ZAzs
9Bticulcy15MrwJlBo2pETmcKkVCJ3mBO0pmTvbMpy7VYme/Bs+GoybnsBbHd5gx
4HflYzRGmZqbNUSAE5neiQjmELYGwHfj9qsAE75OWiq27vZuLyRBmFeNPHmymTtA
UTz1vn0zfqsTwQ2By+MTB85OdR4qg2DIMjaNhEhVqwX6AvU8k9LHetQd3+w7gkGa
funOt1acWNbenXQE2tj8Y6pfZqk/IgH2pctR7IZ1TuonFG8d3pFburCfPzBB10Ev
3WMpWlCE1fpRxeZxB7vqyn5U8B3qs+FV1Y6EpvXzMLxJOFMUlQekGlpyCqd7vVv+
VdeQUFOlVGftfYmw/2EheWShpIvWR2hUa2VBQYAbZFd+CrYvvKQaphFgYKVRZhsg
pTbSEKkDR5EpvVowMIy8Mt+YTMfsmOZdgbYFBbtq4KC/JJL2rGgO0qjYeK3smOqD
zKMprXiNhc4+ney3D97Mw3DtGdUgy10Tbz4a1eZB3hCcF1X4z1FWDkBkGBssx8ba
JS7JAuP+i9LZenma4Fq5JG6gyD5YuOtgEvGECm/BAvRmIP1sBEFTc00YIAS+VRfN
47QccLKJGPL4rrntd8HhtZ9/9nhMMurJn74Mx2OCCS+jIbDf+KNAyqfxqj/6Xivd
reHmG/+svIoSp68sUvaz+dBMFM7mcMmrZ+GxTK7bu/q8UhkB0dH+5Rb0eYhUQ/ri
wR8DFwzafu6o4epYfKKG8GlAv0PuEcptNfC7jqpkIKQnfZdT53wdd7NoNn6HueR9
lTatnm60gBptiTuJFcAY/dgrxypx0lqQyHp3NKiHQkYkWkX8/vanWpIdh+kIFuob
mKC/l+H3rNPZKk+riPfzfrQ7hFBFxmuys5a7chYz8LaZqOIX+T4hfErTzYXGQuEb
Sj9Z+ax0eowy3oo99E8uqB5ojfVsj6t6MZJpwxhulEwYy3F29ec8ZcBJbBHYSeSf
+WImhPTkn6Y8jOd3HBON0lZyw1nF6+yCVYzslATdKDHodaWRwH+hQik1ap588jYs
JTXE900gkBursy8n5dE128JeiSrJ43hDBS5qhV9050h1xBseWq8uXqTC/DJuWY3N
VxPnCsAu5zS/OBcsme/QQKe8eTeGh95Zo5JFDfPLFaIbkk5QQKR9q2FC4n4WYd+/
Zh+A/RwZV1kBD2FQMRNqibGjDAdlcZlJKA9ebFl+JR6/edT0qz35b7OYuPeQ/qeR
VmKjObItXFz1BbP33H1AFG2Pfoyy/wMuBWiz9KthDrmWRyD3Fll6Tu6txdafemPO
WUTU2GF9X469jTw+U1SectsCJHFugJnc40359RQ4bV1e5g/nbN2jLlg0mla2tQ4B
zu4t4k1RkgV/LgxM4p0cy4YcgKzqdDMWE6OdM6NnaBKVoIUMByzbHfxqrts5YzvP
Q5R1yeXYNMRYnRBWJB9iay7LPfwLfN6nOtzkR0I2/5Itm7VncxhQ+UiDXvyEn5XQ
+jsEZUk94GXWocsR9GEdW3JqFFbE/D4u6wdmmMwWlH/ATSfGt+hxPpypd/p7wxEx
xlHnJ/MpXAUby/XLpMzJq39mp9wMqxiJ7izv32LrjMdP/Cvzf9SXg7WKrX0dDR3H
VpvZjW40NO4KZDzWuuX4YtcQlNPcnvuwZkYptiyZl8QWQLv2+wsYxM002Gs3WWBb
T10uHdH/KycAZJBLCqPic1P3JUvQTGjV/Ik2Zy5GbR3/Sr8JSizB/tQyA+E3Z/jQ
Q+IlrC7eNuYdFixv52xBqoJHooDcw9K0oc0jS6CljV9a6OBqxZ18+tlwdzSGeffY
cqFkiQOVgTcPMBO/NxiO2yDQceDkFyqFilx/pqa7ezdN/zfpZvLiWH0E9z4oeiM/
3lfjVlBDsubliVkvraSwYorOk/w4CVy7036XSRbsui4qeMFd6T7h2JTPVr8VdA+e
/7mIk0YdEDZ/ntSlFMAh8o6VCRUfqE00/yobL0p6lhD/a1cLSI9m2nukJcUY3Hos
P986QHLW2grt9fkBzHnp/mWFpL35HqdDu7+ko5lrqoJL4rM+3t/wvmlS+N8Br7pm
mW827msgasbIhNcmxdN+YLLgL5ac0yUDtc0lr+MritYxCSCBw8VhZVodFtiO7dPx
X0LCih0b3gVmmZ7VQ71pkDmMbrFNlDrxHcLWbYUSAJxTKV+u4Mn2o6mCUXIK2eWz
zI/6w5lAwRIX68xbPecfVE4pcUVbU+cIqA3QkSNpDBJuIa/ZgP4XClZ3Y+ZAmL8l
RMJT1NHda0rKZFn3YvCdpHlY1fy7xyDXMBZd2bmhAo/5ydA6rcXUZJnxC76xjkbT
dUdH980uuZOQxxU9aZVS8hxYeC76B/dtXh1BjZvAFfqAiu6ZYcuc/wWG2JmWNGXS
lEnSu2EtXMA3+HIW3v+gMvexPyNlsDb1oDV9RGwcOLuVHQD6dmBBLPO6NBIfMS0M
TeNXxfrmRny2D3JvoYHC9qrv3BerVMayC5hgYaZNejEeLykYJob1cQvuo62tOOPH
TXQmvaFj4b+wMBiP/I/FugLMEB+FseIZK19e/Px6h7bl8wEMVTXbC4R9lyOl2Ob3
zcJC1gQcClQKs6uysExuuDHwZkD+ibXQTRG8eEs4tgPunaLX5lC04vprA5HNmBVh
VRtnJ1I5Er7/Yeu3KiOiBEESsHiHE8+gkwxFFgVaRCgoJz31DUv8+EkaxmDoQjto
0gCROp3oYRjWm/FVj0nhu/3KX1W9dOaKJA6i0LoTBcOylJN8VLYgwJttPhHvHgoh
ra2atlz0ETY/dg12UcOVqHNVf4Zxe1KaOaKlVK11Tzfjr7mOL5kcOpD7Cpw+be4U
yaIs4yTnBjvN1H3f9QKkiJu+oYg2T4mqSu5wSKU8iC9+WeQvN9No/8l8/brkwADA
RvrWmFIy6wMV8pWeAjRuRjnqbek7Qq2rzOw/axn5zZMRmvg/qRSe2hYzHCgrRQJW
OAGybREYaXJxTK/Vph1zuxqHcLOhz7WBZQoMre3VRf113JRTWzB3obwOWDADlXHn
Eue8RrkpeNsUfk7x7/gRooEfKGmrE4SX2dgyd87Bnkd098PGfTUfJQeUY+aQrTKM
fdJkTX558nB7geReFBAw+3DOR5fTlIDMrT1nz5BVa7ak5bli+87xkCOAuj0JOyZh
4DQt47FomYwX4094erc2DcXA1pelV0hVA16NGiJgPQgn6tq8eMvEZsqjMaSWHbBt
wOrhPYIGBdSJsbR/k0fObaHFGJaMluUXh8Gj3ZpBWjXPykNlHAju0+GJIRFW60et
1QfdcgXijaCUI0QV24pFVPHYe6BNreLUOxXsVLSBeCox5LBsSsU4nDCaZtOAHnwB
0dPh7Thl5FY2Cc+Tef9W57WA0HTrJvBAz8kSeKPVGG9pW1Q+g9m35yXuJ5HWoXqi
bUXHz3uytz1FJI+tfgdbNOHBxUBU5sBo6Tw38Xxk7qfY85AMLSBlEbMTiR0itm0Q
mluQlk3zvzGXnLab0EQn9uGi/BY03ZaA9yzAyRy9Fu2hpS06mJlGeJEdTgWPwz7u
/CdmB+aX/B9xlKovBhnd+KoXVXnsF7RRrTCd+QroZXa5VudyejaKTFm76/GS6cap
jJFgw5I+dZtHpDYfdWEsCnjASxj3zNEUSHYKWvB39ZOZXCmfBYEUiTrS8qQtY1WY
0XKpS2P2LB0cBKLjfFsx7KNUsmclRWWyM8FBHnQ/7izAgsGLV+NfOtzOxABQ8WWG
/26DgzWz8nhYmqmJlisnEPXFDK+p6VIcnTnPvhd2rxRm/6S0kGjx5Xp9rZW/adWi
C+PogStvQZ/AImbpClGz/VdWPJUKVfTA7LmB5m1aPRXiYXjRiQbZEI9NGgWTVFHP
qhYlfiaaZ2ImJI8yt6uA0MTLw70PyCqzSh66GE9Dxp9ned1Dcap6b6QPNjg3znGR
I6isENecwvH9rmUqky2BQ9j+dl92Ij/Ns0uvihvGRPZf0IQxIf/SiFxd7BmTAHu9
+Km0rd1CHUuMwb3icf3SyBrXbyTgGhvMl0Lu2f1gdVQ0PeOZH2MdNy4jvGgqc7fX
TC9ZoH3PXdrGP1moOzERCWuBk9HZdjGDA1qRkAUwM0FHIXKGcwu24rShE+GUJ2eu
96LHeaL/D7LTt6lFsVM1aAAQbjev59igGHidoWeekdBakrw2sq+mr+AVFdrE1jy3
KfWnPFpIdvcJY6pK+Hd7nTT/gl0ULCWKnKsJssNYBN65WOWYbJc/kMXcTxPbD9jY
geuNKWoQp3wmxzMR+aSHCmxAN4XsPpNQwYT47IixNirbcfYRWBVLCm1NLkL6vuD/
Zfoa3jNQtKlMPaUTc9c61ye1Q9gCKyipp157sG+lISaJI2zrauoYOuG/txG3yWvU
ZHBkaivgJq/MALMe/eysT9WgTvyZzYuK/fPr1HuqKNq2YC6oTijQYCSF2ovenLD9
XgJ1W5NwcG4fv99XJDHcUKbn5RSEkizprtpo971jAFByAPC3ZjimFNb2TyHij6sJ
zyiLdFTUDEvF2WFVHEAoAuNRqYEsvIJno/2/KAsCghRsTsziInzBGUlZgFkuUwyY
wNswIDQUpma2MfehnRT8mbbFGe8JLxEuH5TxJ5i5V+vJGeem1pahJr3AhS3uuN47
tA+7vQ44l+WM93ucUFBsX9iDveXBWbMlX/42ZTGoAJtdVBwXYZbHhXjhS+AG2OWB
XXzYVg+43y+ATdO8RI4P+6qXHfjtjgO35dqVfsu5tn5gUmX70O7Z52BiEjastFDh
l/+xzSdgiX9Gepqdk4dGntvgqodmSQVUGJtLVORkk4ZdrSP/7an+prhviKRN4GJX
/QjOX5guKQ/1Qaf6eCyXZ3oJplpl7To60BNP3gsOBBy4b87Bq6efSChIKYNFKqBv
9r+parv4zTJI+OBGR+67cEjbs/Lb58TIcdKjOlf2IXXOKbyxxGg/NkhOiODkQN0F
po5RKLqIyAK0+rhRxHStkJsxMgZx4SLmBB4zvEN5VJDdWI+PcnIpzsqbs0KXV9ID
oOUaj+Ut5EKCVTP9WHANDlXIFtoBZ3gu886H/83jrYlpjmldqotY9h3aKgKVXlNP
j6NvG13qEAJoCdik2QsRfITHGsnmJM9wB8TyUnnk9YswLlUK5hqgNI4BzcWvQ5+B
6cADE8RdDB18rpYy+dpfQetGhi9f2vTD7UTz4QNBXwt1xkRTDNDeCNrnd11O982F
nhrLY3g2cHErPjNzTCxRIEbTjvNrXYI/A389GwvhURAj2lG1VjTzEcUtPsAPURdH
GCoDEvNUjqa95twMNq+KcR+97XPCHlUEfp72JjYQA/2oqk50bDfQeeR/9lo5VEO0
5mzzdoKRCPAR565f0Oh9GgKiPJ20IOVWTCHGQIqbVxTSp/UTFU0+ykDZnmb7/Zgf
DWTtcDviNrvR314PdS6OSmowGokrXH/7kBcgVH/+SiIofblAPhtvm4myN3r9NXSE
0IxkRSwh/9oxYJle4+hYpsc7oN10BnPv+fdq72mCPJ3DMtuDW9hBzXd/tapoSDk8
f7yiD4pfk0FDVFAndq7cUJIME//l2Bum6vSBM+OMlNwlWCpKC32HkgXep2yY5Akf
bYxWasqDA/pUOl3HSQb0daH5q5LrTN+JLXFouSZI4xGKXHgCJaDgHt88B43BTOeD
Gy+ebwYxTw44ItwCAxF/2GG8XGOvYzlEU/SWvlOXaxgMPt8Ibw1csS0JogOvH5Ka
0XwTYumzzFQ/N4zeJ9xUtgzeNJQwgkk6d8JJEyCdNZG4HgV2m+nOaD1a1rrfz1E8
iHr0JP29DfGWkQs5CYRBKMlEUNOg6Ff4D30iMsN+1NAs6uwk7Gey3S8RPpAG4YPM
OhFJ6Q9wo6PylsCeE9DoAIjf+PuEsCcbnljRIQ0j465SAJ/aeSPp98cdyaCT2LdH
/D+2EVxFYtNlkJhdGgMiZ7DRIeQIENTgyVpbFZ8WjqtsjWveGplvqP2t4cgpwULv
NOcGXJKqJCBmYSZNfLbNx/NlNjNlwfYBEQdw6RDx97LP2C/oW1mLUN3Ka6L//NfP
H4n6t/Xmp0vnTm6gAUuxbVAYTpm1aaSCiEWHO5sqWiYbJDWpsHVPsyDCgNnwu8j7
e8ab4rHhzvBAJc6Noa4R0s9RZXj0bxSoTiOH3w8KCefmpt8I6h67RxRGYxNnCP4N
+QZ5zEhJk4WOZT+ueBJ2UnZcL3/I2+B4CYyNVbY9Dc6zF6WFXW7B5p68BqUyFVz0
dK4XAbo0aJUuyPmbmEFmQn8lYE4/NrbzKE5bxZhqffU6PfpLZ7JNGw56jlCQBK2N
uxYIoZeV5xf3JEq4zmrXjzviOoIMDN3SmxJXOOeg/Dh5mPWwd2r9HwiWXmzdp/1d
2K5FqWYSZOhY5OHzcYkXelgvHoqR6ZA1RSan+hXHQpnxfPDh8ghX0wF3pe7MQgnd
8rCooVd686+3kMYfCaNvseNlqxwhh2npdDtwg7pMLHujQ9sp6jL8eNhVnIkVHyRT
IX094CdsN0/0OXqCdoxM49j5uDUj/OPsrfPZs0xpKRgOiussbH+eHtJTbpt0Ojla
WIHFDLLaizhH3Mo3RwLGx+7wz+/rUgzIILQ6KErkiPTzcO9ON+KpNqKVSwJDp46I
w7CqLD5LSLVmTTASqvomzo46guSZX0fQpwO7Ge/Gw7XxozGG0YlepAI1c1pcpbO1
W6fmU327EfrKo6Fe9UsLx4e9B4lNCFamQQVFmDjSOUxpJIhzI69nO1Z6AE6QGBl1
UKz+2MkyWOSynXKOwL9ShE/hc8lepLuG8AS15hZqxtNrDCcTS9nJ0GC1Nm9PfKuF
51p3PeT5vxxBJEA/hXTBwvzwflEnSC0+kblN4S8w6zZcPXqr0SalBE4f2Id/ZHg+
SpXimbcMsCm0nE8zoX4Ge6QSqIAc8svE6NvVsDTgMSEFQOByBK5TYxSfN7lt+KsN
ENwy3ZAfVdK7Jg8dQwPHEiK+e0/tMw/djbIgFa92YQw+GU90yTu4PbZsUUWa50de
wpmYmX3+UHETCRBGssP4Sp4z5jAU2SwjfcDOYoJfrICEhQcd0Jy+5fXywEc2YuYp
OeTqDFaegErc/a1DNQYJSCIb1ujm8+igBZ6jmXFER49xQHvv4maOdeaz8Stdd0qF
bdlv0uiuokpuP5KcSd3bbBjwDtCWsEeRQGtNGQ6swV2Vra/YJeFLXG8IXq3n+roQ
2585GTTNw1Zt0vzDfL6fWRgKi+AO4F+Rm8CBZzD92b3nKMBc3teXA31v4zh4VMwL
Kmb7Dt7EC49JQrA2khqJMGHClqdjElusVAB5qOCe2/e79Su2dy1CF7n1Ohwv6qaW
PS1t9bJduRVO9A8HDVaOq29X07Pv3jFEiJTKR4GAtn9IXj688/r8x55Qh34fKJ1E
DnHoe9LRV6ytGW8IC0aCQOIitQqEFu86CmhWwyYSkla6fxf6M6I9i0QyD2dLmY0Z
3oFP+EEOE9kfvRndagmU+b9tSGLQK6IFfPeEXwvszNrclo3948o/Ai+4goi4BnJ7
H+xj0jtBEkeMr+mGUc6CN0lmEZU1HRYYzkvc33nuhrzZkZPrH7hVLWkiZjUhN7ff
NEmqXSFdfgWpU12rOQYbr9qj974alLLfkXifDxFT28e4DsOHpKiujXy9dxsK81vp
Wmbt84jm4DjZLCN5SQOJE7AtJfuH31TzcCk4hUtY2aDFGM/Y1emcAIjwIc3d5/9T
Cp5HWfHOmCsDxPJeWL/XQapd1hGrZFl9GEfxTDAR7Z/aa4hZKi/n/06p+LMY6RrX
S8PkgoUJpE/N3xo80L3nkSek3Y2lj6qeDFpS+8xhGaC6IbFmiXgV4LRvfxgSta2R
57G6FsQepzbB8AfAgoDwvQcLg5dcF0ikReSYDdvLg3QLxk+MJIMQH064Mg9MYQ6U
fXp717XIxz+FNgttYlb9R5bb1z3HcNDt4lTSp9kPZbxixTD1Ni+SkeXVCAaHKcz2
eQQknVUwD9H9t89PFQso5SZ4jE/z0+7oBvQ6fIQJF53kVkCe6+Y8IkxhdgmN9Zyt
SoWKRZzd8H4leaPlU3IqwP3rmZY0MIi6Urn3E6VqEVCOqSGIYA3fxX491m0b2CsX
EnGWpsLCiiNaXKENkCwuyR05n07lNZ+3Ql128BN31f6JKWY7Kbj2SZYFQNlvCr9I
83R7ey6XQlpCunaMYEuqET3RjkT5jsg6BU0LUjKVxn3B48NiaQaxPWbA3SMw5wHB
IExYkWMwZ/UoUTAuv+Lr4UYNh0gqKMnPtD59pC6/Dsdy8BYa79pwjA7/pniZJa07
L75v0iFkm1oYKpnDqphuUFS9t2OV9xKh57IShGipksBLwSUIZ2rY2z50o5UBv2P2
MbeBnjLonOvrjroVijEHXMZIHpX0q/WBaa+E9lE6gCHiQhGRdowK3Klj2NADZZ7w
7gwRTqHmI3BE6HkfUlr1UDtZ8nEu+SDKztq8c1hcZm20OF0c33651Hks+khR6IKR
yllUPPmVXKFIdioCyxYmtQOtIlVAe6l7ilbhN6vJnQ4xNs+cpSNC9Mcig6/Le5em
GzCEyzU5syarYT/hfSRhJUH2x+TyxjVLKm93dNyLgyWohZffKR/zyVu5i0kz7d06
zexzyWbsa3AoGgJNU0NDenDaL60sXoLvmp+p/Pn8/8uqU1OWqoobtBI2C4KIQplq
AIKfDPs1shF7gATFydD0y1xW2INhIPflgILafoO/l1ymyTNrVgyBCjHzVpkyAtfY
8QsO8jx7JwM14gVd7pTULyJAUYCpHeDVEsdBp3X83ypZEyQKZCdFZ/Xb1e6Q9OyA
2xwBghBCLyAM3gCEOtkKVzxkbp7zmc0oqe6MqICkrK1IwroA8NxE3pNvlXirbQrU
GQVWyIIdZmJesyVwEcqYQtHiDYPHhbsCX2oMf0Db27ABuBHtbSfBKgfjvjAh4P/9
l5zcpkXvfGx5H1OE8h4DzKqkoyfmHgX8n2dyvrsId7T73sEbF5FZl16Xklqqh7d+
jXl32f6cquh4Apir/2Sa3Fki7hXYdugtyi3pRIXctgvrV+vNwBxwcZ2qYl6rFBD9
5IqccCBK7fZNPCY2G8nCkzlpDv8DWskdtIQ8LLuns0+qgpp/4uvZ8G+QVe53MCeq
B665C4RfQA0oUkWFXuSGposlOt3ZSvFSEIfpQM87AgeP3ZvgRg+ayQ9uaDM0RGSC
kmtfXZ87pW9w67JQ25Q06sOVJo/DICnxruehffPa9K/SO1AHkUMMnrFbhXWucfLi
hq7/Avwm8T0wZSl6jvUkilOTJBNMGt/lnw4ZNnpMfR2nrR48gd7hEOy8KWYABH4b
9uu3GOEHA3sgstHdQEVWXS8taj4M7ZDE+qEsE55+cP7YjWg2seWCqFB2V83xo0Mb
DnMLoRpQkGm7cJD1661KsuFpnuB5zhmYLa6T/F3VRzAayUjgQyq3zD9fkukoHTqk
+wI2aYmZ4JOWUSFqzMFnO6rTmXLnMdex06NbK5mQwVt0XfLOGymotA/28+iBL8v7
f8HRgGac7E6XhqM8qNQ4pO+2VIUEe/heOYmdeo/Q8S6g8gQtwkwbxZdYLMPuXkFK
IyL/1HwAemd8BxuNNcgu7b6grNmxoH4JiQOd5IEKF0xXFfkYtHMTf6d8JKd4eAHC
Tx7BD/o/MbxxwZd+UP5P+z5M6ukOiY6uH7VEqsdt3keUoUzgCS03WRrcny1von/w
WXu9EgP2hRCMrsd+DGiQiDMVFSuNiyesZ1tqMRY++CIaYCiW8SjEoKH33PQyLXVL
VIvn4z20FJzHicVM9eyQ2pw5CzLmd7/8m1Z/XyIjwbREBEwHOwrqYeFS9UGejzwj
hRbZ0mJj4tSiryssKtCwQK4KY3uOKkWpdHWung/TGWIp19KsMpcZ3IE8ygrb3Edv
bhTh2y0aOgFh5Mz5ujKHQDlhOrH/+0Nm5CagOtLt61BhNAIG+Co6ySuQAJWqlXjv
daDzal8MJdCnzDK3wXOGwVNYxtJAZ54SiYr1GEGLxhF4cosH7R73ye0esQRff1qc
xDhjckVr39dxErLznPLjtBbCaf90CXRfRd/3Dmhi2E4e3/ideHIChqPqjYtOr8EM
4bxgn780SQKUQvHB+HnMXsYWNejJCCjHINTCfDT/fDRBJDw2enKUSWp6gsttb8fA
ZuzqJOI3IEh9aBG7HXwnslHHPJdNaJVt1+gpQFIyC1aNpOYVlrgbqEgwfbg7S1cf
+guFU3QdUHXJTDn99qi18X6NtVhhgocyVfLsy29cR/Ah2LPOPhC8oWJkN666wE/u
xRcYib2Ac/X1dvQOPEP+vP0pZ+GCY8W9o3O8CmsJAnDSC1wA4EZplQp2ZC3BQvIZ
2zRGQcr+dcmQk8/NplbdE5xV1hsiDaiG/1iPfizB5z0bWoPirr5vPHeVGwx+if4n
C+BXTdVpxYu4XblcXDDArnH4cjw13F2brMnST98aEV8l1eC5wZmEsY1Zl4J3MDKX
Kw8iElKg1kBsFlMzhmyt81NVnRWYuFjiZv+dswIu/IMTIPBagr1v8CxHtfPedH2O
QtSJLSSYpd/uDrvgJNVqCtXEpieofF9dRK4PUByAMuIgB8F71AzJgNI78piNvwlb
nOAHyz9HlWfE3pSzZw+GGGrTvMXV3v000DqqtM3kdlwkGcphPBL5Iqc+xRiTyuHn
YoQt0EBY6i0mRA70eKadV5G9T9Jq1lUSmDEvVcbKpETG/StQZhaWVE/xdh+0/lTi
aZoVQwweyQ54LYdXP7DaFAPZvN9Jrgl2UszpicJiOFos/XW5UW7NgEj5PTQW92+D
F99ILYCg06TIDz2tFn3glHnGSLRA/pi9JMusVnrybdXSlYj0BkotyD9u7DB/KNUT
MkvMrzA7b1MVkFMaGrOdWyfyjg2O0V2MvbPVvqEdYcXxv6PgJSPQf1xXbj85EX2Y
cs4gyHPL9DeIdOrfRuAvxfRh/Tw37BfT6up3ROM1QJquUC8Oy67qbt1ajDfoM7nx
bic+1PY+nPT/soljNuHDVNbWLkwtE+uDK6GwYHxPGIFY6ikNYOy/YqItLfP6l2eb
Jm96dw5MeX5D1xccjcEISauTcVCMWjD/rlTABqBJU4b0eulSm6IzfN9jzPc4e/fJ
DEfEhZpMa/HHmInWD7GdO9bT2578pfN5QibtnRoKNyzkVjUQxSGVXp62QWUyrrd0
l87ymoOHxQGAWh+O9NzAhsuH+tl5rZ/TJoL34Waz0GmXOsqsX3+G9s4RinaJzdSB
nNHA1CdSNL1wHUjcCsqzxrKmNq7OSZ7y4hNkPCp98ymnQSYGTd2MtJNZmbcl9ZQy
oRH28DKkXqyqy4IBIC7k/5HR+DdAqpmCXd3h+wqxghGX6zGud9SSupNsgo4HzYVp
lYBbmkQQG2weE39l9JM+wy4x14PcOF+DZcBw6TAK/rui8SEbMp1C9cRltqOZJ361
w2DY8C4mhgD5OAvZuQYzEe61J8/XRNRu1Y6Dx/VMUH6e+2tQhye4IUA9fNovmue3
0g3l7FGHeFhzo1SnXlXuwncDBhHFPIu9WAnQkjaqVhUUgLj2BwqL4imHBstlOgWb
ZsvUoNVBLu/QCgog8m3vcglUB1Sr0zoKFZN0zHeICLlGhLWE0mV/iFRZc81rsYVs
lixK9bpwFz3XPuVnTMyrAbkeqyAKojF9DDfCWd1l7NdqblshLzmN/8imG3OuM6SY
Q/nLxeIRSNjNyj9Qirq6X4GT8xaVKzNVr6vMq8GSusUUjJqTGSGTI05SRNbarv52
DxqkWMU6QyaOSBML0BR8BE2nvR22Zhvtb1o9q2CIh1gDpbEHdqLo97QXCFBiqnxp
62VzO5mIAc1z8TC431+JKpcavlXUmQ3Ob1VOIuHEVu7ihspIe5rTPLFJNXT/DrQs
tM+FRBGQ9cs17XPR/vfcx5xLGeolyQv/z5iRGjDb6WmO3/M2Y4s88+uejA+RGfUW
SWFd/AdvznnD3XTFR3Vo6pXbMU0cl4K0hmBhPAeYj48jndqOCx7HQKV3kF3T2OrJ
hcnyxGcBh3Q8SEITUboPN5MrecS2IjRdM2DV34PkXTgKDV4lgAzPczS3Qs0UfqBC
qbI2zi0MkGk+2CKjZ2BAg5jtWbk7NZWBzPM0n6EapWprJlPdvP10ph/2FHwYplRb
GGnokinutB1O7tzCBlVwwns2xxrTA9jZxSQvwSS6YQomceTZsO5HiEryAsLvSBQg
uhQLt79nBRgfPQLqhA9BhwxvK/X2GrmGezSfabWD9e3wRcwc8Nvwijor7sKwd7kq
P1BQhP5FCmDSAu/8+itAGgdtSg27IY9+JyF7VmVcqEeIyMhh7XpKwqt/ltRcIvHd
2QeRCNM9/A9242U/bXKNzo/9rhLOSaJdOvdDWQTz9iNiIPudj9QPsOwVGCYL8ipm
PfcSwkbhQjDWZIQq3LRKY5TeJhRNow/sI1f0ptOiIq+ZFXlXonau0GovcWjLO1sz
Ap2+4ena+eJBuH5axPosbmogCITF/qXZEp+Vd+XzBWUXsx4Qz1uCRZPb81CQdtDZ
C1QJntxaH7+dPB3+fKRPNepet45mpli+Q2nRhY5KroZKC1UdAwBgN5W889XzEtye
sVlP33kUv86lxDMKudDsaAjMNqrBbYr6r4XdcMMaqTClnNolUtwRhD6G64vuEKM2
prRqzpgrGg8b/EkM31VRWf6s9N9JNevQoS54nM0TKVyH82MjqOXy7k5G2Xo2OvMK
9onS2url6LKfTOnm7mR4NllAL3PiHqFvZiVCX6v5jCavwG0jGxw9FT60wkeDQZXs
Hej1esafPBEv1R0/sw2fB5bDML5PWp23rx/P/qzh0cmF+GgB99mPzwMUihUvHqX4
k4tRfZ+4rUygKOi2tFWFC1siq21mFeHEJNclr+6eDwvlX0vRES7YnGTw/iJ/1eWu
3lNzZwiv4Bdtt+zOjvJlxX0/VAB5FBnrEeTs8zTyNhOTXVqp4r0NgmACxrqfcnqt
tCFgv9rM/YtMrZY5jXhPSUKw4w97BS4XlNTjZU1Lo9Q31eBFNaGM7a4S6CFjaJZu
OUtsnQgEs3XACX02JYzyZB4JRa9kYrWmenzXRy5UX1VWYWmhMqQZjqnhSfgw8Laj
i+8fPGJt+yjk+mY8940WJTWpcSNgLexezYGZVAMwjm94ha6sX33q7u1kC1VSgq8b
4OdX+omCEYIUGY4xTqY3GbzpuIA7l0m2iB/ks01vvyM+R7pJyMeZ6G8v3tw98JzD
cPe8oA1NV70g8UtCzQz1+G2DKOQMaRqvw7E8n85AZFKdnysT5sPkCizjmuCY/3+t
yqioz87WrA1rcidMtpELRSxveb/zrgefLSTpiNVsDvTqNtS1/DumPwXTEkCKP53K
y0yyXjgdBvWxIc4kGpyNDeyBpHtd7HRkgX5VdDluDZEo638Yr/8l68PlzXapAY4S
j3DyXvSMC/mdyo0pbiXfVyWCzlKSxvw6JJXMLuYxivsQTQpSwx8iXhmVNHVZelpI
AVnn8eSptNSZVZEoAiZOngXld5NaUFZa1Z0MEYFpZsvhsIG53VQXoKV3rjEW7Rac
UAYTiPyqVhs0j/7XTDUApqq72lyv/VpfMwkDkGvU519G1G9fnU+V0nBRnrVPwMOh
RyKZ/9fGGy9ZJlHsPxHYi+313/CT8v+TPipxAs88LW9CNZ74t2XNp9PZjZiP2WJa
q1IbJhRlE4jl/SGzdHmX/v6yjFtVolS5AsVJbQVnvkj69sD+p2g+35fl7+jH92jX
0KTrz9gEY4FUPWodwziX7U/CdDZghSvbdwr6svbNHTiOD57DyV83D6sxJe0GG+zW
ah6LJQ2AxFNTA9qbamOpK2dfU3KkQmYM2nreYKQfeK5ofyephA6IJXEGUeHFVsvY
UpMEFGl5keBmv7nI5bZSPjpqy3iabd1Zfw1NKotuRL/uHFwP8r8vFaEu2QdZnxgE
r7nd6LDhsJ7pcSriNj2pp2uzWh3OzFhH1iCGsPKyQGHiQvl5AsIiHueE41lWtgcr
HKQ/8IYGHML7DA0vi497c85gUOQ9YzS5wFZ3JCjIbc1HilzuQntnQ9fJnAJZ0cYt
XZYkmt8uQWwL5jilwflFw8BTkTzgeNH2MMFhH0EOSzHHOhrrfbdrVdv/F/ikczpD
7gFsTt2k9W3ByuTiXn2DrjS6W4GeV1+kJAuCSDoY1Hv/Te4wlhM6ccl42LZZKJYz
2KkI3eIYwJ6Hec7gyHb8CPr/DCQGPAqM5Y+SfsdI+U2bEUTFZvikWBOBw+JHVRjm
iYxVhfVXhQTjOIPX2+J2c6ZdvXnAoADNrR56oc2pjgw8OQu/6AQh6dn1w1+IcKil
Yqbav1Cy0J8pQ3t5GY04TSZQ1L4NXgcSN4R7MN3fA1KQOiUjaJdAyMIQPFP2fVKe
q43pG4tBfDqmLxQ4eyyTq/jUt9tTzAGxc9aaElmKS8LNm1bNO8wBcrQakRzG6opI
dsOGKjX4qTcIsC0QOaVPm64UXDLfzfWRl4UsE7Umw8zYv2kScLEURC9io84mP/1E
2uSNjFzvOwXSHmvuSNUibDszsId4DB2dhTw83br0Me76TDtOd+fKUP1gXAxzetFe
SGNwOX8slafk7e4qV9MHNB+6/Z7etUW2riZIZ3WeARJ5NXP7v09gxnZ/Sr287s1E
bJj7obKDBcwnN0Xb5KH0uMPq2KcL7qc18WPWEHKMD1rAvHb6d7SOdlrNR7rwOvuv
M2cP8sC3rCn0bClhcNi7xSX1N2Px8jEUPUMZm3h1vrhvbEddJk/D9QAzZ05V5itX
j5nAfBVayrF721jzTTlmqlWBnOnahDByhs/TR/pBeE/wdZAAC6Tukt2vjsJIVXNh
/cgTiTWTRNpu90VqU44eBQgf91ZrPrkQxsUttrGAiiKpLyvIdkpElyuXtcLIik+a
MbtlLBJhuDi6TfkdTd0WU/FUyXER6fNntJQQTQkceDx80GaqBQzE5ehZ4fOqOO1x
1qBBRfaG+TM6yl1ONsTg8QkkHryCz/LvsVxhiJCo+kwYFuCwa8KxDQRhfahWC6Sy
DXqXH797z0PxGKbD7D+myM8xCjfo3I+h/SC9iYEWfuKmvpzNoIzvwhgQ3D/QApgf
YQlh+dbzPkR9QW0UZck4gydqQma/vbbChGIpOWSmzd2QfLHqNrPiofgpcj93E/FX
AXUJU+GQp1O6RQ4qX1o3YatOpKpLD8Y4XtmUgJdSHpppJaQNSKkHrqBMqISVyTE5
3pVA6B1rq8HbcV8wP2Y5PFwXyfWUU1iZCnMAkeNadbCCR3fG3aOdr9cIQM9W1Uef
jk645mGjvaZeXELj0d+PiIzoQfukgAxnZaRQo4sae6yEy5R8VxtGb3EONMHRpJuD
SA6pXn0LbRvdgaXs+Dry2p3DPfvzfZ0O+21rSNBAItqy2UOysA6r+UxaCf0E3FDm
WT48fwEISp41hBeEH/50rlvd4NN9CjWzqTMBG1GX1TO7jIeonuX5kHJw5noHHx9O
XUG9/7ZR+Kck7WhKvgpb9RpW/XaVGe48U7Tf/0tzSdKTs+2cT8pT7L/QsTXrcSWe
2/jc8eOgMKTDN2/O7nkflWJMZZHUKegJFx71AjK3NB9UHk6RBqT84todwZ4EYGaM
NJsKuOORAe1ScTYSLVWI4er20jEWPTQRl5MWkCmP5MpXfiOwd7VSkrJSC5/PNUjl
+oiGPOHdv2h9WuNnRwGUtnvdF13LiC3bBNPMfBrtxtGve8/bjkRy3oHqsOR3t5EG
MXRfAiqhrWEQVFbCFs2HSx7MOLxhR85bEbh5jblWWR0+thLwokN2D3lOJyhhjmm6
kslHiJrMeFUlilI/t/Thm6Lb0fd3aq5w+wBvBe94mNU8fongMUgeJLcY0qd+TGxG
wqTDTb1aF04AH+5yCyu6WFklA0VAA9oVJqFIAY8mNaZonYIISQd2sZaBFaaChnXt
kS7eZdUr6fwrpT9gSwbbEftkrgoMw+Ry0VaeodC6Jad8eMF7nWJP/k6UP/cqpkHs
uVYoiehwFGhrWj9WkIsyrXK4ntSgZbCUMZED2VO6bDWEHcVLiVTzCv8n2xgu+II1
UOvNTGzj2iy+joRP1nJe/68FlvRRz1zeIrORpUnbg4AbpSQ4VQKSmIxC63ELHwoy
9m+DGjOhoJ5XJritZ2PJABc8WxlYviimmehnyDh5eLm+SsAqgQ4gKPR2aDPLAqaL
XpeCsWunhcGaJVU99Cyog7i0XL/AgTIrhgvygaKKVlgpq/KR+6Z0SJa0OTYY1F7W
rRNOoh+XVCPd0PKmLIZnci6pw+VQPDVuJSL+JrTdxjUyvREYe54MwzEiCQVrTIv/
HQ2POIH/gg6mmu9ai7wm4PWVAR126npZCnuSl6+Fv34kTo+nUjJYhGzQpWKM+1MW
w57MYi4Tca2HYT4q99hftILgMlL2ZlDitqvglSJkHLunIlUPIgTCjm0htY0FZVhC
3fmU140N78xNd2Gi2XbmjcP8uImjHqmKQLtJ8HnvlQ7nBwSJoMHhjzuG8bOav/Nq
48dX3McetiquIhwgHOcfqu38hJ/jvr+DfrtEY86eLUm3UjqH5a9vMolam6iOHnok
1ghl1dof0jISS1mf12OZMAJF14vxHq2VQ0FUef/EVW10jwOUMJl1la/jxmR47LAS
7zuRiW5LQbzeS2IMYN1sk0F0Hc7tguBL8RvKSlitTCZxCO6788e9+C2cO3d6Xu0C
XLr8doFjvH+D0uUvZs1xss+aagpnTSXCOzoLmPzIAI65e0dBbFjPqRkDmaz65p3W
0ysbgelHpDH8ZtXs9/0NmP2D6dYpqXxCnrk9GxANCKO7xA9O20n4yH/YQWuBR0gA
I2LJPnA0YwJ9jNjvOFZkNdRBhXkJxkpEHw+omBkP1KYWVUmC2UqQrpp5D0Waux9F
GnN9SealYTdgMF9ZH6v4mb0UCac1WoFebiRpIWJJ5cUNRkbdOgMZdGwZHnzww3N6
AyVwDPS9c02eVXKqeCJzKbw488jy66lk+6GNB5DuWX88n7C5goRvaDAU8besPLvn
cPSwhTAhhKZvl3AZ1rwPlZ9Y2f1SfnklqTPyz7bzV0Z9qZHP3EO0QvqbNtCMkyWM
98hbSzwHAkVVGvoHpCJWHakDrAIZZtpBxXfu9YcbXRV3oF1GzQEJ8DvuEGPpLqRs
p9ytCqTAVDX8c7PIr7gN4/mGoLu3hVi8TuHJ9sD5B+5af1nNBaKSm79YVEiY4uzZ
z5Tm6ByilbYhKWzyeS1Pl2hJSNZnWw8W2CqN4ze10jYD5mReR2w5QOmKQjignjqv
f5le4xK4Ywr/3E2wSYcT3EZxPLk3swblHkP9Lroa66ZSuzyRkIQwAppNg+LEt/Bn
n3R/tRmE4+KbWRcyybdqWbVSwY4BEhYkOAQyTdaDtLJB7WFCOd/SSziYc4KcltLV
BEVdR3NqBBWxlJe5a/7e9iJDOB9pwNNly56ljGPPUTfzzUKYUjRtwLZDKNdEWcWo
h0GEUqzO00PpNOisoXRI8rzMORTB7vMvVwCzSNkl0Ik42nOp3r0/GzsmsEzf0oK1
2Efzs8gs2IRZE9qQTexfilgH7X3Xg6LT8d8EPLoQU7iFT7E3lHMTBnINp8aF9ZHM
eW44/Djwcs/ujW/VTOEeGrIBLLF2wHTRk3PcPIuTJ3VtVXb5KKRmuAhiT6WI/xP+
NdObFDZYas4C2xOomkksb6z8fGfUanwWlWEdS32jifsYY4LjQnVy1MJ7qXushMAP
IF6lY6bS3m2PbFXiW+NdRIpzlNgp1h8TBfmDWXVqQoxXdb03epZx8rieKxYyL/ZZ
OwZ4MkVoAdK4/6ccRdPLuxVCKcjViNlpyCpwpoXRWNCGcusWp5iuEZcVsKzm6T/A
IaQc2MRM1Wt0+2m8es0QN+rgpeWU7CcqubkYffVhQW2VBUGZc/HHdpF0UQXBUr6H
C79COoWaukXY2L9wcWsyCA5AOspXIu+uhiPn7VW94tIOvW54PTJm5a9ENiy/A7zT
m6Gm2GJOOq2r8nrWtHRvJ009LbwdxcgPO6cN5nWZZFBQmGeLPKcR0rG+4S75p8S2
+JPLfSRcoSWpYmhUSb8TsWY2GJtola35l9vO6Pu0i3/Dk/geYIS2Xl4N9YydFYQJ
vONS6ypdbTL8IE/ABHgJ+J64vq+QDI1f9YuVaBxeoVYylVas2q4DRfQm7u6rN+yG
KCcAt0VPK1xLcJlDWvwRupUPAKRFLYI/XJ27PpBRfnRsJfSUy1NMgFsqNbOKRpaU
RRnyQHMvPhSPcx0gb83JpbdhqgB2ntNT5eoCl70UC3VFrSjIjHlGcBGkkYzNPPdu
uajQsIP6TjsgcVT04SyR5Nvcu7nGbfpjy8fwJ4XMJgC9EBsfRkQ1FrdN9st4p97F
pG/ncVSiIGmW+bUn1VjJcclHv7q4KLmZ8Ogdg/MFizFyLJ+Prj0SX5JirV+vvy3p
qlbgY4X1a6YHantPGlZomLLfiuaQeYNZKdNHhyzOEuGaGbGw1bCS7pDPTgp3FSiy
Sy7OS57hvdLOK6+ensj18arAyqEKFHOi0ySMmdLbI/7HdYoHcT3jW2rEdAgOn73E
PzU9rKHt89t2cIe9rv7x/mDF+Bx8SPVdlRq0dEPtIpslLckL7knxYL/clHCyezhf
Fq/uEOWe/q/Ojbg3lSuAHtMX7DN52PihHRHryTkMvwVUVI8Vf2IsxjtvhSsuvS0e
ALTc4zu0Ivm5Ftjv342gO4br30ovdh2JtpvNt1CLI8dW/z0au4UhsbzWijF8fFFy
mdQAUUNLx3n7wvjXi8YHBjd15Fkbx17hiPrI7P6Mqej1mH/MpHFJyZQvP7DhEEFd
eP4li2TzXQy2zH6y58tpelzBxk1CnzzlTuEz73xqb+T3NWKbD/+7pQVkUgvNg5s/
/yIg2m6F89V+VtZayul09lE8yNWysMmuI/o42ouAQi12ZVX/9XDdBx4HChBl0VJN
g9AEXzO+JgTZ95kNKAV9G8zmkB+FJOnYnIL4pUewmY++vzJA9h9xfNGh20rurSg8
RXTH7Xg0o8vQvekPPYx4qMZU1PdIV4dzCB9Ep3JcQkowA0Ya3aeo3loGkgkfKtcl
TWdK4xC3AOyiPmIiqEhVujIvMffgeoM16kuxdKZU+ZMzYiettS7iRLDqinl9pYaJ
jQHE7ZEnRy6eQKR0/4EDaMIGJqK1sh6fdRMPKn0I740Sz0gYrAB2Nj1sA6cb9+qB
Wfsn6WB79Mh3rKi6j2gmzHNJDyNX9O7r3BB/BX8yM1rCA08IIzQ4YXCeTGLV9gnY
LPZ9KMa8l3ew24s2+U1ZoPXSG+EOJWIyhHKKHDdgDbgvwBYHjWf93RA6d3TJiPiX
s44Nm/tcguEWk1wYpqfn8t9uiyAtpJKWkI8oBh+1M0r5i4YKnTFLFNklImMI2wO2
xN+OSR/G8hAAWg3VnJ/OGlwOlKCzTDe9HFHCLn953+rdlMT1IhIIC2mVqxANFpPF
CZCQhiHn8flbFLIVTR6xFj4Dlu77Wbc9eI8i9NHOmaebsjUktMrQQP3rPtWyg8SY
V9P8NSoGuArMpU6Yj//rYNmLbZqMueQf0SymB4zuDQ/6BLO21mbOLoPqFna5xL31
SnSOfWJs9KW5T97G21p8TfqVJMxT8qC1mk7bi3zx1bdT6+LguKexuOR+iWcc2Cju
NnAXWGHbzikjFDx6Z99kJ49m2WnezS96xsPvv4tBRKpKq9+mN0YeL7nagxyMHnte
SLv/4WfhSdd7fAp2oVythTzmbcQln/PukBrbwH2K7dywYVAO/SfzX2lV6L/zKkk/
LgAFSfq8GxNuWaAWCujSbGsI6Ip4KoJbpO8IgybvZwA0q3ooHVCy0K3uNKfB984x
E1a4zY1dq6V0mk1qezph6Jtecy6aSBrcoZ1IfCmSo3R13g3coug4w/b1FnYH4k7c
xfwmlNTfJtVr6Cl7MMhdFmYuuLvQvwP4ZTbf4VCo4dBTAXhj8l9ennWunW9hH93b
dTGvhtBa+2KCPkWFWH5eJh+DHvxsH71rwvrZBvvC8prQZ0JiRRP4xSlvg0Eb3i0e
R4YQKNXs1r5J4VsQaoF2jag+6mxUgXX4ktWIpHoUNyyy6XcyX6dFczcGAIKDuzDm
b6iPDnmM/j2nyk52xUhQRJK4PKnSaR7Fru8KLJvGVQqJTz0DXVj/remY83lpxa/4
QpcHOlSFLYFy8qF32oGypFMMu3qqv/pO/1pALS5fKRpjDZYkZdTvOCUy3xzG/4rR
7RNT7DUh/oIWwAJ8iuZ8oL21eYXpcViSlV0YJwppFphWQpKeChd8vy3yC/+qlxHf
eaSOGcmXHFs8APUgTMFS2Hi4/AK7stWY/aGh0F5AjVfC8nRa1CwOY55cNyraFIDe
EQs6FmBVmTDKSOY+3Mq+cXNBm4+bZQ1l2DL4CLSmZFRTuU2rE+IVL8cuai8rSy/d
/XmjP6QPJaIlApAwRPPwizGc1jKnvxM4Zi1AC/4K1j2Afo/CbZT4lYn4VuVKmOn4
mf3yoiQHNImSITOhpsQT898042j0EsIr4hz6qU9T1GJ5oVfZiw7W8pXE2H6tcxLZ
nCEeJLCiHu/q6mh+pN/BiCbjON5DH81aP2DjuyDOwVV/X11732IcmdzS/8LHwtBq
Fi2WJUcRInO3mzcsxG0zI30gDFB6quHkO/tdl0vOKdgB92g7V0zP6LTdF39EcXjH
Z5wYO24q5sYZYkzQhyKK54SHPAArmTYkYyRsuh1HuXOUR6ed3ChfrGMCi2ZWri/V
oX7/3JgY2ghM5KHTi62lBDaNlwYwG6FJojCk4ydxrzV7zfwdwYbCA6ZOt35m3Vge
blVa0y8uDwiawsZVmmPa/GaMjl5dAtZxHXW1NzhDKxnOVi8avY2SXxVuH0BRQT3Q
3lxxGLrGz0oHhIQG1ZeqmYcTcaIrclIT390jPV1OR9awK/bK5bdKb56G8B/vR8x7
266RUn3ZQVpJOyp+AG2saHM4TbcA68NfKqPxmtT4jzyJf8T0mA7o7mSJNJ5AShd5
TJUPdqieZPQLnwwM0d2ybsRtppP7xl6FZFl1TP1wNyoPyB2IH6x6j+4yxsW5ThiX
tyOwLTnhhAdGaqaAbN1v4/strJQ/VRR5/0SrUU4QUlPXFpwWAwXSmtH9LwH0gIdO
09PLb+hf6tF3xY3SMvEMiS0qNjdKqcAy+sGVZYNS3YPWSWMT3LuCdTFSZyi2UuFi
Rext+2dvhQEQI7cBewe56AF1sJqkxUyK+qkyBzL2WIJpN3U6NLpv36OCdIdmW1GL
FruY7erLtisFk9x5KE+3oO7EhJFJB7To2ute4kfEJEEBPLgkrp5Nf9zynzBlUrJ5
mryDgUXeDX2DnAVPDtH+gbRBGFYCc5wzvZfCvv6gxEblJMF/gLBREwHtGgPh0mi3
4V9Wpnk299+zHIrgTLNa0A3LvA8bpIoKigbaOVoCjNxU3Kn3UppnTLD79LJ2SVyh
pm6vemn8pExBv7eQ2S8H9rtmg/vzvSsnx4VnQqv5kY7UlzWP37zKWBkRHwPZt98H
mLsiGne/z2fUmCTHfsamqX+Cl1b5NasXlSoujPwEaX9sgXRJAMSTLA9KokUgDJ8R
THU+/sHyDil7FYdSGfGWur6RckYuQtDQG3Et2h9/iYtS5sLTRRG7uhJmuKCcdXSn
iKkRPqfhaIca0Y2UEVrmSmPdhd0cAYhajPROiiMjuewGjPYvcTFeZ3h/Lx/FzCgg
GAenNhSpfASsG1xj8SpArnE8+gMNiSkgugG4Eee4p+e4cuU9X3Tqbs8XW5CEwQDy
3bXW5A4eS6Yii/1KV/l+9UFfDzM7WC3w5EjdjWVtArpr4p6/d0RHdveS2tGfVIP0
xDT2OcI9ia77EVo4vQ8IvpeCb6Kd2AvHyip0A1OH9lFKVG59G0kYd9C+5edTYPli
XdL1Tf8+XACJzhA4KHoS7XEX3sD+Y4M6eZpirjWZQghMNLU+85s+v6i7ljUJqGDm
S+v5MN4mDPShAtq7E1k5fbo6jN8ngqjbeGJBOo0OR3FxSTNa4eF4ejTHuyAa2/p7
VxA8Jh57O0UVYjInrNWs/DxEV7cd42HxeADqDgqYmKsBGHaIlQjCKQhMhCZRIL+0
uJbfCw0/q84pOC/qpZn+sJa24TRDUzCjoefAP1qhscOjP9WH6zhOl6JcW7zTke7o
09Va+OG1TQRFARE8RMrHy2sgoy9BoK2+6NGpNjgYcJPZNfx1K8xML6WhN7Hjmb8c
1tIGl7q4rpHBI3Hrvpt0c/qiaMQ7VfLOdzLYou9QvlpN1jOVb5T7m7w6/Qxw9UKd
wv5a45v9v3ZNMdO8M2TKdrayQph1tPA8zrpGVHsO6K4TNzxhxChb8lHDQU1ne3/J
wY+Qkj7oq3v57JgyZMzQVbVL7K1J6To8aAuWlIEGiLb9nG/xTQ0E83imtldmbZ1t
tATF+LpB5bQLjZrrn+h7qF/IZ8hhEbLZyZAGtYk+0mzcchQoBdZTFi/ytRgBK2uQ
UUyWRip+2emjOOLRy5rTOzsI9bPajHLdnXLEtRg/8lSJj/hX59/ndlrmhGtugCSO
iRajK1PpZ0PRr2p4L1CMMVQgF0Vjn51CoWIp/87rByEU2z0R8L2oUv/SxDdS6rn1
cfeAmig+dXVeE0L5GiYbJH/nc7S9WXTX60/oUtdsoFznOwtcIJOcflG1mi7O/gyC
uHcJAA2tJnk12wfbNleeP9Y2bSOfG/EEuvtYyFrepDrYp/2WI4am0V/NzRNdzR8S
svlumxtemoLaFWvxS9DO1fhAsqdbcsmtdLuB/WR7PwSU05p1jRsOvJ6dTWdihjif
ZVv6ufwLCwkx+FJLrMohr37CdMjMWJmp3gp0L8kwO1nhntgdVsTr8pxoITlXK5eg
trr/2dv77EsGccOgMFoc8MCGrcQDvfL/qMGrh6E/Zc/3wzbj3QBhluF2kBBqIyCq
RoF3QQPK4TeknEpYS7d4+BoLBwLMFTqMmfQerKYQ6nnFKpJXN/uuxho9J9/UAvLr
HXguUtEzYHWTafWJhB3wRjFdxm96QuC8hbho8Wv8wnehtySg1pItEBe8K5WDHRYT
MMp0s3/ECVWkSqtYd480i4mwDpgHAjM2K2Y5QGWoYEmaPcqZCrXRJ90ae9IWH1mE
eKe2efl5Iobdr3h0DxfbG0MynPCvVLxU9BYPrxG4JmOa4OAzA5Cke+7fhWXX8ShZ
cD8fA/1PR0sAsl/BjzOhq8V+B5BXI0rmmdSxrjJBfr++EqiwgZ5DlPQLUrNd1m8n
SjdZJEBLM3812jJNnHv8EHlaxLTQzwbQhBhJYPToHVfa8CwJ0tfFhuVK4pKjbYNR
y9XDRmheJQBaQfEdWP680vRM/kKqWnlQOL9qvn22Szl6f8NE3lOujbiOiteinMUj
OFHywne7yEgecnNBN2o5KVuYjovaENKFmmwVrw16Ygyngt2AiarDnYPTwuXqkJFf
QEDr1TEZCPQyx6pCaNYCLZ/tJRVkE0DkJSGoCshR3/tvsYzt795nEO8O8b+/czJW
eNVwJuU+tTYxJOc2eaRAVF1xoLVdSB/4KQiUFRISyVoEpv0SQkO8gBFgo3PVkIat
tKyx7YLDPtjkvk5ouBxDJ8zDvSJjqlKw0QQcOfmxct0f0kxXR64A6E0YO8p/eiBh
ZxKw3QD1hrKFC2IpXJ4U6JYOIbJ+OK1kCo16/mX4D1QG7xLflseJCB37INqg+Mi5
5am7wtVn4C6fEHNZvz2OldaY7LaDGXDHPBrGuZ1zSwVdF5pZNYl4hhwkqxElQsiQ
zRyJwPc16bvONo31O4VD8TSjnbZxQ9gwmTQj+9w0fuK8aFmUYoVkEbR06afCCnv1
eEWuJ8H4Qp3uzmYPMDNmp3eURK6zcV8fOnihb7qJ31ZyToxMO+I4s6Cv+R4E31PO
owD+qNd27u9FRb+a0a5nW6ARYNd6LRWE5lP5TbRH96Lz3GnXtUAbaT7ilv3qVbFz
/DFxLwxQ8XgNlGJHbYaAXGuakuR4qXHxK/biz9GdiJbybXci3Z6uhluQwJxzihfl
2fS+ZvV5ne+qyani9+4r/qz7QuOiFht7MykDC8hH0GCMPcMa+1rFztHKTcS+4HP2
WJHI2x5R+KcPgUXsC+4xyIwbygQdzS1H538VGzVMOci1OBx/aqs4spjviC+1vPvY
H6DijKJlwtcvkjbxMroksROQ9AQcgQkrXs45zedc3TfDbt+vFQ5ZcSnUlimVqMXx
3/9UpdiBiMp2vPd5/zJVKgZgxuIjkmhbjPoIjfM634Xy08LQDgsoYsiianOQA0eD
o8JsYWjUAdlMJ4oCA9OJZO+a5HThTDLmF7ngAKLVycOyaQpgycDhkDHdpNhksDOy
IIFLKGqN7DySldk9zZIYkFpT1Agn666OysTRDxZ3YqsrIkz+w5j1ttGio+Uj2CmU
8xhXAFaoqFQ92+4GOjoHv/0Qb5tr44sZHQvDkT321adpLr5GEipmZGJXfEirf9OD
VUTu1HBX+OPaQrOpqEHTjZnBFdjkhCRkzDLU3cwp0XWpKO6/8v832tRPQ1OqJaHN
ppx4cvdCP2HETpBfNYnUuqWDbKgirAN6VEDRV2LjavoGfutD65W0ly9EK0Zl6+2i
6TVFLK9mBYokProstD+Xj0P2b4QcRuaqQPmf7bTVhrk3C/FlKbqiwI+4YyLpWrGh
UF5fPLX2lV0TFEPjH0cx6AjMDPSptu9q7e2sa7wCO1Rz0EHjy0+alxweBK+eG0qc
yF6JfjhV2gQX9FDmnQTiYwa/aOWUWA+vBUClfmNOiX+k0ExmHkJMyre90aMmQ2tX
WEb5W5wmrq+FxKhAJB3dpqNrAftdhfqmJ/coIk+LLRKkTcxPiS8jPAjOIWhV2Pva
JIP3QlODXrPpSmtsLXXeURkXn+kuz2sWRl/J1m+kQvUD13WwUSkL92sddyl3pEr1
aj1KaPXkhpY3HYsTv+XVP3/NLCjb/Zm2yebxqU3Zq/Jr22QGF58JhAE9c+qssENk
me53TrX7dEfnUBQbGY+2vRVXmuPXckDr7MdZQ4x3OOMkjCrYc1bSRWFzar+Otyd6
PQOfywqvzFUpspX+b7iRmYST7At/PQ47ZhZ1rgcM85P83gVkEMCqaI3l1PWNE5XL
m/SKwMQfYSGbvGEGOdpfafKJ/SmChDP226SGy8M8nyYPiNWqkvRKwlOiUpQhgouI
bI5iy9cSc42ab9v349XdpmSmCRA8j8oj1hb2eGzupZT3gS1IdFvJOw2gDLmSOzxw
LlHU8VPD72EOlmyu+WXe2QDEmss1Nbz9kQUY2wfF4dEaEwZcRC+s4wreWyq1lJuw
GPRPA9DfpvDqfeXLerZTF+7Jm/It/Xwg72Zwa1MUDsVqstlXLgZr6hupkmp49e4R
P2RrS2B406lVVxD7enVXZPOlaBvOO/wLCfw4ZfZgWsNQHJdG7SXSjPqnZ1kBYRqT
obsmK/Mojxk3jeGEm1CC9Orvq77J0I89Djtq+f1+cVs2qiTkwjM3DFTzMUZbldls
chzzSFiQx0PDbKwH9AFXi+3L0wrzHkSix8/lKVKFkpEgw42p7sJdaPiY/fh+yzL2
zP3lvUqRm9zNpWc9xwEhjKybxpFn6wdceyVv6WZhAQXzDZ8LchHo8mKHzDj4+69V
6Vj6PjCUhNIkXO4QeZwkxK0M/7hvkRAg+cJbmeLYwKSWFo/OQj6pi/q+p9n4QlIA
eLlKor9rVxdmLv+/oXsO0bjLkqCGuNxVEWxiG8yUan9y+P7Layk1XwFTN52rgh3e
uEi6BOi56Ef60Q0CdL/MWwRUa4JXVFJvdLbzCezh+lw1Fqjt3A+R7H5E7NOmHaXo
+nie041OlXVxMikTnNK/yzd0Y7P2R7UyRjUKn6+Ux3BU0hd9uQbILCWzPqppl0BK
h4SjaoGirL8mjaUbSxoMpdtv2atu3FLk4jYdu9VK06NKaQ69fKKg6HPvoTf+OmJf
0NPPD6//bBDlc33+3gGOqYM3mf9nYp7rRt+eJ9NL4mTF/0xE1SUg6EAiK1U6aFec
qAPmFWxpgztCWAuW9qRuHrmMoPLR0cz2HiTb91Fr2GHlt6wYkOf2Ca2Hae0E+uBY
jM0J2fgJ+tSaCdGweyz4kx0hwnuPnLgxvYGo95KlpeTqj1q+8Pm4aXW/cmlwRTNX
XAq/vupmtU5iLNzSrp3bmEcory7M63FNI7L5AnPPKFriwOdOnp2kqo7FF6i8EQ6n
q3uLNDCIPETR8Hwef46swZhpvvpx1LAP7jgFkCjto8mj1qJ9X50Hwi/suoh87y/L
6HLlFrLs75LnlegyqrpguBq48eOx4Jc7W2ObeaiZhEYpjh70rpyxsaefi6tdilES
vJ7El818qXI7cNNHyyf7xqIDjCfZbNPm6I1EDleqydf1hJ/L0bOFNKUY1Zez6Hx9
L3hNXYU0OaxqsglxEJAHLay5WXHL0sbjiBUaYJX34ZUqtseYSYZW7cugXzPdSFLs
D9ALVIYl5CkWE/NgVobcznYHbQM4jOt5vzfpK6vfN+coFYHPp6HdajchVZGJIKUm
Xvs7vJq+o+wZozbjZj8e5QnNSJeEpx0x3SHyrb1eIv3Ldbzba8CecNYJB5iOcIJn
q/3S+2mpW/Af2k/EgGyw71iJqRL4PdcOat3hG8Oy91BMp0hbewKgOSlaNmfRHrj0
MjOuqC7xz0wsb/kLBomgjj7gjORQFMfW2bRqa2HbQa9pQCGzzn1w1UMAzAM6pc0g
2L0XJ+Nn601YKFmcTV/I6F8pNXeYs6y8IzDjH4/pbELpdTSyT2SKg9IXiRArvhw4
1m2c0VCQMouDXxegxUFoij0BaLrz7Ju3XRJPrdM+XEUOUjCtGO4sRKKznWfG0eDM
4vb0Nyv9BeFOksKCiV/hwKU0TbTvvRqfOqg90xBX+Ffvv3zLp+B/lZoVYWAUW1Ew
+cm4PMSK0KGqGGrw024CWzzfYu8Xa1svov+EFGRIxf+LoALzqarWANVPcsDqAgKZ
Qqm8BUVLNpnWXrEvpg7pQ6wcDAQa990bWui59ZNqaiovPeagtm1SruS/MX7F5fZv
d3g1cQRhaaspt+11zdSSPSfXXs1ZA/cCv6/h+Bv+xV2aX5jy0ALrAeef/4dOn11U
utuZGikvzjvWvfgPUwq8cDYVP0VZERKlg3ymSGsulorazqi4vqxcmBzHnYxFNZHb
S/im1J1TzWCi9hRMgLu0cI16LE3nZYVPLvzqEpupk2dPMresp2roLD+cOMwBKjRL
Qdwi8jLcrTRJsNOl/JbIZ//n7h79a0vbEPb8x9PBUY11Hl2EXr8vIhULyptka/Dz
akunX8IiQteCFcPBwpxi+kDg9volc/QYUx3G5jHeh8Yb5LV1DYs6Xbfm3tBpIux/
Ohm4PNLIwRoyAeDYpnCT3bhG1aFzpCGC9Lb9yQaHRRWpFeTrNOXuDl33ZqHOQu3/
aoQIt+N5M0ld4mO2A4RW1E80neIt4C3Rd86fmvNBLLyEMSPar0i7i6ocmTDy/Qut
+spRbOKGqYZouLsBMC5dm/lRE2a2nI9ogw/66eMwvd0zVwwSNHFSgo3XZObF5qMW
AhKoJQlCeQJOoWb2dXnDv7HmAzUP5Ma+8k6UjWZ8GrX8Aq9O5sJFhjI2cc0nt6At
/D/ePHIcfpsI95MIUol/35/XkbPXX2Z6tOZCr4JvMpE4s/UABtjKKbsNxvvi5fPv
TXs7U1CqZhCVjrZqUbAXl5npcNSsi0UbQAUw9af89FYVbi32f5OXAj7XZNWj0Ed8
IlwPfyeY2oIYATdUGyLzmRcbeiif7XTcdmEQZiMUTkS+UL0W4hUkeCYLTRbgfb+T
h+B7DALOYcZ1Rrw9mScQdqgexQYcRDsKyXfHv4JWsL/G7FASOkUVqLRZWACrYja3
kilZaO2zbgQVIc80ZDni0DRdiVSvTK7epdvP0CVaBWcBpHhLe6viORGHydwCJBs9
KLagjCZutu/thKZnUnnFPK6fAQqYcQukXZmfhML+zTTAa/AFhEDdxT7TQoXWtp/Y
GPVQfnr/EmeFWm7Nqe8jAxqQIMj1aw1muPESXPykXUvpSb3rCuqWpHutg08kbZ4y
eObtJbbFoRgBd6PuCKktOw3jjIi2jbL+u5BIKiCoXdxx9UDbhuhhyen/KX1zQgDB
y0yOJIbrSUKxqWUqQaUudyLFx3gYJ7+/LHCy7NbnvBSJvPbJGqXlgLG1+9Sf/25X
xIuG/1lYNReAO2xfIEWfnpCilcw7ZD39y5yycyKSajNCoYFxKMcZ01oSiroPoaiP
RpN5w46aNQd9YeIZi+j9Xh569sTNYOHSIKd1vJkRY9kBbj1io5F7XvvsFt5LLxPg
H6jb3tPfUxgSjkcT7+DNj3RCkiWUUMTo6voYaJT3XXdmiDFoBSihTc+0FB0iDiJ1
P2Sa75L96/Aoo1sRNDWF1mQVYmg2iPUwiu6Qh6S5A56aEoTx9+U54Y5Rlu13JfzJ
RIOrduOyRGnSSK7bhyxhyuULnAPmEvbCoyw1wG3TVHCKNNGunmx+fWIODYQBJ5Q0
eed73UsJQIvSyu0otdsRFdDKxhDbo/BdHnuHkUZnEShDpbOarxQgCOpbHB7NbGNK
i8wvqfimSa29+d2Qo0OJfP/cpfDBuZs1DU7uFDNLq4we4gMdXYy1SPQoUSDV4d81
gAhnwCthd0xgh14MQ47TPc0h08maCGqTQJ2oQPDzKNQVcBOGsjH2sSnhCj2nJcVP
4ITQgjvqbAYJeoJjDV1zWUugPp71ehWi1Jf/VMPUfq/DE/bON8RNXQDJd3v035KN
E9Co6vjcTlglg579pYJVd/5SFCVJ0n3TN6F2kc/W0IwCYo/31/c0c0DObyDnQeQj
+paGNlpzuFqp/lywI3Bz3iR7jju2jLScZwQ/DFL5cERTT9TzXVvc8Tm07kkXyA5i
VKiySUuB6H8LVZA9jsI1ytCG+jmu26A+evSSjlCL7x4pttQ2nbBEY4ZLWZmIwndi
554kuiKq2fWIdo3z/vpdyc7byHmWOu9bA9InjU4zGgVO1yS0j2dkuTE0JRyGzDGM
A6+y8iP9Vi4QqblZOxZiGXCusBN+NPcR2o9BTZegxrK1ZVzVeHRE7XzncFHPokb4
K6Z21YIdIl9du15LGuu3rhxLUjSICcpPZrYRJi7M6shBoAVFUWZCn/9ux+PRsk5j
0hGTaZ6Rn+oVd9BTrBSLnlPE5RFHA510ss0rWuy7DUXgR5/uSc+MXLKsB13FoILh
zckMEmphCGNWIX9MAlA+i3vRh2Ibk5ovCGDtYGXAftrO1ilFF/ec9X5zdvJoR75v
Clkp9DIbTXkvCscUSwGmpKI6fxYgSz4h/aPle1Dzqtc375epf2Wii9AhgzdYGSiU
WWqdr0qZgExxVnhcuk0eQjwzmd7isduuk9a4p7ZNfcht29l+rUDld09N4+hQFnlp
KZ22COW9Rma59tKZ7mn5lLSUzKczr6cYd1pFNCDfSRLZ9hrmSv8nI5EsFF/ao4+h
x0zCF2+T1234ef8nIkpOKdrbu9OvZu7xs5S4gO8KWe19ulvenyEOxdCxieQzCkIj
bX2rtmU3NeolRu5I9WC7oJHGm8TppdPehr/R1gSHN3tD2DDBTRCBtIFePNIEztHO
ysJKYZVPoHeJjaze0bi40LINXIkufNJxz05OQczP9ncwZweZpTEsKHdaDALON8fR
mZUg5uR/rkZE2gkomQRkHwqFZZMbPLvZbVuBBSwiK+fLp/AoWVZbvVJcuWThxl+v
NoKCyeDJ6kG+/Ci3abWpNauRzi9C6YzI2/SZ7RhXcBLSKx7RkclLDr5g27+kMaTT
NYdv/Z5PEnT5q+Pf/SjflYHxQKuSULbm0PITAGm+ZJxZY6bSF/+95XvdiSWYRtSU
aUlvCxfilg+Jsj1Fap36UH0tVvFSoyvQ/HFfNTebMyJXhBc0LdzxFOPTrnUHMZ7z
VFOwY4t8KnXwMSB8Mxn8NeYVe2m3Zm+kcn8ghOS8sBGwwNl2Oz4mLFLoPU6kIcWB
gvS2dMvGNSdAG3YdKm4l8p6U25DT/xhsarmB9E/ocxsQuglBtNeBmAYBVp+N7T/z
1keb9RJb6Vshzek3W95SQAmsvoHZrv/Y3lD0HMSTI5BH+mg8be2ogYebBxjQwy9A
aPmmGHNVLJ9UjoxYs+WKdB3LsOwaMPqq3L0NNiwZu6/s3mXYP/fJZ6eaZ9KQgN7O
+jFpeyondAGTiDMeNm8xTzOJUYCa/dcmHhoQ/aphI2V0aFNmf5jMrVHCkI7ONF+4
s1XRvAtE0hsU6/omUcbvnVZc5ogkJJthgwZ2tfPgS4+KzAQSprJ2chsblSWLAWu1
R1LFNuFoaGGu/BujqBzueYqOEHFJKw4B3NLKjPvvl41EwOVDy3rff1dSf6U5Idh3
mBAfDuJN0VljwJ2XWXJWgkKOxA/KNC5P64KdAhzHG+mZgyxyz52JPazLWVF2AM5p
jyxwItqhRNEn6kbF1NTeK09AHzIwGsNJfJz6fdxu0RUcpxQBw6/i721bqqtK6TSr
QIYlHUYUV/nWUhJ3OdJGlxJ/v0auQHLrxOKBA01sfCIyyGkzuF0vFqzsodRXzoTi
5Nv01CBKpUjzk+yAl5w2AmfH8Bff1zJYDPnVZQ5mMuB8TkvlRmjCamXJXCP9r6rZ
BdgDj/C6PCf39t/Gsl5IM3u+Eb+duVTI3bgc3aa1XC/+v7vdbAh068LqCNOlcZ/x
miQ8Yao6Ws3TSqiVtFD+SY4K8FipUuZZwYRSDm636UH01mJjJzWxOXcYz+O7lx7k
c6+73s160KbaPzZPIIK+s13R5bsI2v9PlX9b/Z2nRbiNBl64nlc/w1ds1RhEQb54
E/VG1ld3GrPGllJH0pmvEcUqipMEu1OzkAUYDYv88VOFKkv/gF6mlzzOSAwP+fhE
5ZdQC3mq8H/JL8dkJtIq7VatyvMGKi0Fp1VXciOoQsVAIK/CmydAL73jwGKGHfgm
N25zLhD6RSOJvPCkT6QT/OipgK9cPH9JkZKHWO6Qr//8sIx4z1cxKzOWuVmP//3j
925k3kHCYNivMa1gsXK0DACdTXyEKI+kAzILCAmL1vVdgV72mph3O9wbAJbxLLMV
r0Kk3jzsob47ODKR+wNTKB8kM0S3g0etOZxc1hI+gvPxxholJHl9wZ3/Qc0IJXMn
E6RRMgdxesrv3puZymOMYY5Kh6jcN7fyv2jXiP04/aFmHbs4zu49YEowivNV482S
mlqGcy5L5vHpRKNQFe/Du7R6UuKqx8S56Hz83DG4LYKb9ni/kLwTKBOgJeoc1kq4
A+PSATh+aIIMbPUuzO44L72cuyx9ykKqcM8TQZOjJPa0hMkk9VkmSWs47+UeyO0f
2uk5nhbg7uzVgGHAcj3psW6ePK6CEMQpreKKZURsu34tKsCzp4R7dJcfTVUxUzG4
Nv644+3zDnkGwrtiM3dOu8mPMdYNcGYja634tTsEkNcDEpO159/mRMKBeJNkZWtC
NGTNVR3ubviHor5cbCCx4PlQN5ALWA61fTybXKdSxHcZu7F0aH5lHY5TpFoIY+9z
ZjlAstAURYELKA6JclbLS9zfPyx+25mqAr2LOO3QrXvyTHCKOtS8TYlp0nQ1iZ65
0MJ4kIK3uKP2N0ZpZiOU1Ru99ObAPrhxX9LolQqGqgwIcENHPQDhqXr5b9/vyb3u
mqyEXofb4gNM9SVI6EsbfYHF6fGo3kja9KsFes75dHy42xO8yAIbnSgTuVhmq0E5
mJYv9qC15j56LtZ3gYalpgYhFGrwFRR/6uqc7FPIUyXjych6MTIxX/W1gVnLXh46
Nc36WbGXJLqAJyNRCFD2/LggNcMNVVNH+iWD6ByzFCOznZ3IWwEVSnEGLU9r1jX4
UCfiCPe/+x/wxTYsgijd64rqADjNNJdP7NvwC8tRKKn2iCNRu242YF/gDcfuOTpJ
Gr8tNgDX+bYy2K+Cht0oXEuNCzbdqxRGE711EhimrR9IZLzz1bo3OS1sxdITfZhc
pk443rUPMph+ppT1mZy1+Ih1Cc1n0jbSNBK+PigXUwq0Q/r2jIZhyQNlvmJvQIbu
8iwX36eJ1s3RWH37Fzzity9JpfFVR5lcGpV43qLRRD/Hq15v1nTr41sOnNaB8iTP
HSo9IKc+WIdST5y+2a8vwJCzlBk/Q0x2oXii1wD2lDSwVvBvhaanJTqAFG1eUXAD
p7mXCi7GzQ3XXkAE+xKnxhQbx4hwsyrYohgVzlRb1L8L5gNW9xdthyIKCxhCXJO1
QCeS7i3t4oWL8skNBTzYgEKy6vsxEyh5JsrqsulguRkekLLwFb6WziSr3GwMSCmB
JJNtKaepYFNsLl9Dcgl/5VJfDt7mWZVADN7l7MxqAc8p8QMdpMjzU2U17aRsYNF2
miVITZQInEajeyqtOLvB2jGN67vFJIOcGeVGGkHao1C27Wv/bbRDDkUqtoogy45k
e8nlO8GopPXaHy+KWeoTq98ysj08Ks4YVb5PzmI0toI1OEqbwyVtGAZ7vvAghO/l
HmpM2bDgaSiuusevy18bk/O0K2IsOc9JbWmTw6/pZ9lL4RUSZOEUTPFyl4WitB8C
DStk2NASfzs83bJDDYpbTWJ9FTw8smBjvJ6h+k0DdjXfRCdF+6Z0Lv0uLZhd7Dyg
5uW05rTU7tDVKKOxCyGVufsYBQ7+W2GZMPLzUUk0RtT454BHzamb6MbQC5/9x2B8
x4mQV6Lm1M9DrVe3/xadYGjyfzkRLQWVMd8zj1FgqoFjxzI+JiYnBcYo8HQ2YsPM
U1j7LHk+BfaOGn5CeUeXskCrNVt6uI6uJ+eUDRBnqR4bxxslJwTeSX3sksQGFQwP
nOLtuuF7wlWbZeol2ESbq7SsYeMpCdW7Le47z4daesvK1iuVwoUT6YnRdrojF9tf
PsBKqD+E/dTXzt1lkd0MTti113Yd6ZWmt2uguRaZT2sDXfh9ZNwCEXCm3L10NxFA
953Zu/OpVx4MbvuJ7pBkwAlWDwMLVM7H7y34OdO5RpHMdIKapM2sVyIOTg+lYFxX
Jw0euNDzfrg8hhYm1zJo1bR06i/Yr2tyvFFUDiQsGAMbGZWCOf8z6Lhy04AAwnPp
yG3wUazP+kElVoKrQuEld4lN3o1SF/SvUcSlRivFIn2GplTSWu9vUBJ6BuDyfgfL
JB8hBWwKBXP1m5KH3V9gfaWc4w6E7zqLnFcqu3zhKfoOpaW3N69pFSvvjzEglLhs
+oV5jHxjUq5qXdc7c/fLgKqd1m/1iu1IRcadNZO9vEbe03DkjUg/hB/xznSh9j97
gTKEAejorRObKZNaKEeigzvWTaUEY6c5mdXZUAK6pjZWLViO/tG3I4jZKStiBWAD
/x2HLqhKbMqL50DwAFY8jlBCK03DcyUzuZJs5+ALPcnJEVlCIbSlV32o8CQBAv2r
/Q4oa2hCt/jV0yL3g3GsMjMvQhFaa+WoT0huIhjxgRW63nYuOsmgOf1FTxzMHICZ
iJJYPQufLFT6g3mSKFmphpvpndWUJSB94UFc8D7qulEdmdqV3GUVd1GdYPy9euHv
AvIIw5CZBt9wLiSt9Ly+6Q+K/1Msm/FRYmGsD8T8DBvhhKS7IkNbJjCj/Kr9yC+A
e3nm/laLiHxfoO2qPFJzYaAFUKenLLINFOXCTLQpz8XGVGYznStFAgz8rWDNjCig
gFVRNbJfIbLDOnpVO97BjWwOJeveEDcuo0QcwOfRNzRGHY+qJxnD0nemMS5taXSJ
mdkFigEZKimE2h1t0/nFlyy+7heYPr5fOa1ae17j2C3pZsnn1Dt834HQebXZirv6
W4TqmyOspbTKWxycRc2CJlI82ga4UMv9MsDoqvvjE5znqJLiz/8Dzmw4UtgKd8yt
vSVxQRW3zp5JgRZl7CpdmSpZir9SDLXExZJEvforgR++zNpwNj2OAi4ekv+K7pm8
ycydiNEWi3qpCX9Y77MxfT+VeclkNFeHpLR6ZltnjFxQ9wN29UPwMVM2NCbKO4AS
mmDqF3gfwpLcE8SXe86OPhY1g3PAP1V10CxsrBPaTSoPU66gLw6z44w9V/oWcAST
e//6PW68HW9Af+9iK3cOtjCFF6tzYGAIZAANRugHs9XzaYBeqKSriz6yW+eWQNcS
47qQskQyWWZodHAShBGkEUASVQZJmFWxd/+q/AIevZAOz+wBRwZtmLSY1NZsefax
LvqtiB4bprqN0yX/EYNKjJs/st8e5NEmIKvHl9sS53lS6FumHmpXxzTP4lkQEWk6
56myVrhfwZ1YXx7McPAGuxH8afukY0prMniCULn+e71DSOamfzjbh2b2kKp91lh7
10kGwLbo1+t11GkmlXVQpC7gfff+8j5SK0M51JePnFqNbduTnRZG824P3Eee/oQL
4JRTkzDXEBqU+Dgq962Y3jLGfwyk3yn02CxuVhtsedCLBsAnLbAmsqyLWhn96AWu
9K60X2R84PylgdLuHGZ9Gy1FDKI2oqWXKWLqoN2BVih9xHEJ5K1JCXEtR/PxJJMr
RGS9xvNncm1ZeWEu1t5KOgEdU3VEREx+IzK53WumNJuhzynp7s+6WjKT6rGRd+eL
LbR9kkBJ/xlMZ8fKRXnjH+zt5taplV4WM8vWQ2AZgTI4Ou20gIAiraMQmAA7ZlBV
+ZEtCbi3cBizCVbSzWGtGOyGhGbnX8KmG86aLXwzYuXLSWOsHmnFCUV1v+t/VHG3
pM6FXoM6aGz/Oyfwp41i3O/Ie42EF38Iomv3DVL7b5zFBcUwYfUudqCadp9epc8U
5sDma/ULEa6BQnFVWYWDNWj783+PK2VwDbqHyMHeHS5J2r9xqtmcc+3gq6/tvvSs
W2oJtEP9LxZiw0Nafsoi61TR0OraeYjXNTouGms3HnumZ/l+VhnCe05ji3Hpn3NY
sZHHuD1Lz8OsoovtaHDeS0uQjl/Z/R5NiouLsd43PanUAVle28Iw6yWHaqR8V6Ox
GhLFo08Lp/1cMFR1QcRMhGiI+sXGQLeYuB2tqMeagD+7rWOi3DqEMp0OEPgWrWkW
6mPolY4s35E4qT1P6bjs2uyZLXlqONjUDcVzQBsnKgCMDX8qT3v5z2/KgPxF2e6D
+3rtrgOeI8inwjjXnq6ykWsr9fGl0XsQ6lNn54Mzu9OW7nPa+6KyDKmhwVuWLAh5
ZPxIr1cYbjjlOAnndQYHi8kx36/k+LxHFOM8N2ZiuKg2HVA22bL+6kPw9fOdmKqZ
TVSdMKZY6D4sBK/1gQ52vUw/GABS+pIFcl6r8hxRoW4Cc8TpME4oFp8UAdm+YFSx
ZgA+7Ry0KTF3zJR2si/GJp6xmRZGit/0RAhFvrMF2YVpRRyDHJLhKKXO+W5bFfcq
R6YBy2+8Q3+oZH07U2rolhNUUId6dwIMzRsWj8Yohxh6sFC8xTG/umACVNmt+0YS
cBGjZHpwUTNqqSrh1aQE9KztOH6q0/wUzj79aTF3EsZ4L9RVXM+sIfmOnEkH8SeL
lGFhZb3+u4qk5r8TYFQHN43PemugHgGHzO8gBeKFuX0LmFpAwe8TqOY8N+5aBf71
Vj4LuMfzxiQwQeBVjLW9LmHQXokZFayMErhJVh6WAr/OoTBPKL1ZhMeWz3ndSpw9
FHetfVl6rQ6WuWsGT+E36K1NQnGVxGqhCWllmKkgRTMo+wQP1KxLdXFlOIuOqgbB
ZqqgoXE/MJaTdgGpxw4hH0Wmw4rlZAA61rF5X2bXHKEZ+h+VpchMY2E2nfOY7jdD
oemsA0roOugwf+BjBpImCzIBL+LIe4fDkWl4lSpOr1Q9S/BqNc0kW+sgYAEDeOb7
MQWRKZr8mOSNdfWmc1TbNsUVzN00E60X9wAdyai7QdtU9S1sc209xNehxiaDwEn+
yrdlvJr1Ry+IhapK64l+EDKardbYfrV3NMC8vLMwjw8DGejWPX2GYLOOvD8CKbN/
E6KaBeNs39yc9+j15x7QSXDq253wMwQDLMJYntR34fCsMw9Voupz1DVxMEENg3I/
a2A7nNTKfGtahAK1/yOjpnlZwqXR32QtRP9gfGXWsspomlvfulvMAiZXov86OVEy
aG1OWUE1GyZzgn8De7mJXjBkzihH5S/Na7uWdC/Kjrc58MGQ3tZN1Pld7SKxpDV+
CwwWjkeMdlxy+nZwe0WqEAQAxAyxrMqkGadcUY/j2nk13T6bPFyG6JCGRNMBmAb4
SScw7P7I0eJdUmxy/g5qsy7MjnkZhyfPnMuFwlWcCbKBXazSn8kvHX5ONptR47lP
RVzQwHwiftQuHdpFzlpIJfeyl13EvApQ1Q4ALcLIVynRKtLHvd77C0O5QXaWdclT
8SxFkmgUdsEOSjZvQRFKPqZj2V2f4n07qJ73xoKob3O9mIaBTFFK/DD48Xo6IBgQ
ucwHvFCiBO8c7yzj/RC89vx+TpgUBkKu5lIp/mP+dMYjVLXK8mN/pp1afpnraXjq
eVr2E9eQJBQraCDM5dO7HPDPIqbtjciSZ+bj7RbXOuW/d/0QlE2FOX+ykD10bfZR
uy8N24SdRufS61WB1Ho9OlUtwum/sNv1Nbml/v0hs1qXRnUQbu7yP8a07rXAVZrc
ZQzVJhld31nEPpIVj3qIwo/FrDmvZ4+g2T2VLLo4zpj8d/C051vSQcPONldyaxBX
ttKRyKgFVY/094Tz1Wsu8l5BPP5wYHc3+HMh7byWyOj2scsXTQsB2tzemAEyxQ1l
ytuGtxkIpjdVF0gcbmah4Tjjbd3koJeyyftojhxhaVJRnqK+Saj6uemjQ7y5CRDS
tZ1+ZTwzwCCGxJ/ACkFqqXXOgBB+YtKkCeobPXvb3UyvBtHpeb3rmhs5o1yp9YT+
l27avc5ABq5l0RBLge20S3XgUiDlNYltulZjDuNfP2EVEUVBhaNF/7lZklZwGDsM
wmcuuDFjUmGp+nrio5XvaIdk3b9WxRiAZWHUYQyUV8KuA49ymjnbsA0j5yLH9avp
rFPtFs2DsQhbhjLksuwZY4MxEep118C58xpiGhDI/3Mu6HzdlJ+/UyPm2Fqfq8LD
+sA0MxMYLYoGdFopwR2NEBSuHZ0nYhj88soFsDLLahSjAyl5OFFiIvamf5a4gKfh
VRrQYJCr5PquYd9it9ir2Hhg6kjuKx2jTKM4LTQx7EdeTpZ7K9cLwlGQPwxtpebo
FCjEubqXFPKIuhutEZqhpyAGGRuTJXQIQXi0/3jv1P4Vme0SF4OIPFT8WxrO5FEO
aa2XdYTIepCDAX7BFCy2L9Bl01JYcY9LAikfx/LDTNdN1y+Wm4mVqbyue9ja7WFB
+odDNepBIEjhjswjHV9tK5qx8RH+OGROH9am6Ys61txfBGHMap46vDYUaW5BIzBm
PvrrF/jBvAtCb79+b+jMG+2LvUdyahp57Xg6fZaeV+HSVms+qR3lbCWgysv23KhN
NIqUKIXrghgCphcNxnMEwZUjQP7Cnyxd7xXHTrk9E08eK5PU6TuZS8DJP2PLTGoN
gQsTBf2Bwwoa6q8fM/dJ97eRU40mHJmOkz++9HZnBc+67avVhyNprD5bxz6rnAb0
/ajs3mErVXZV/M2Lo/qX+VuHpB/jSWHTNJW6RDTNvqQeBfJKVf06N+WFKl/Zjwiw
jSgfnZwh33qO7Hh916Fv5YuXKccZUgeSw42CNZDgocCtnCArQMomZmDbQbRSvyrT
rtn8ZiCbux6+OzFHD46CICHxxZPGo/GXWCtU+7CtH7yFWL5ACfX2uFHtge+7/emA
3sQA2sCjv3qZpv5q0m/Kx2uNoKM/cEARCmvJRp+7cqNbdIwxcjCFuOCtQsIIMvoy
idUdDmSB1OTsJzBtXzILnaebJeLyNDBu+YJEpobJk7Y5fQE0ypsTdDMHyzhld6bl
n79qEUbiaqUTT/XWD6wKrCLcS76uZvqgu0dtOK0IOKhmo/ojMUfUs0krXRlOuvZX
f/RDtrE+bub+D7kRkrhcmwMfAZAlA42437e19yrsPbEi8PESQolUjfbV5ExLFClg
KmwaxexkTAJTb/Dhe18nJuUIyYxkTxdM1wWz4orBbCugb5QCc0wnqfjA/7O/eaM8
e8ZBtR/hFnjjnq7Ssy/X/LbRX1zxqyBA0miHju6eHwJ3b5Fw6K1xHk/Bks5untvX
Ii55NmgFYUSMDa/kaQc22/za/4DdafA+2Rq6biUqoOHjuRouaXoWn6WtYUEppE3d
jNVchaKtiMRqLeGLiEu6HniYn9yah4Q/HyfLNn2Yf57TD8SGtO7KSNT4oPzWSJbh
mkd8FQLztQYJhJ2sJqQzzBBvBGfMsfwTvzuzT+sknM3lDSam+mkFQ8WggMrWNq0Q
yC8hbtFwnY0n2mmxaqhpVXCgGo2TTiZvgz3o09V4kxbr1rJPASIh1WxW4FnZ8CMt
GhUlMn1ce20zr6QsuZjGAk+z8S+YYvDCnxhp/W6lQ+2y9wYKlitqkV3WmsevZc2j
bygbXjtOyPR75YEjON/BuXjqZqkD/T2BjE+/X3bRhILE1TjXt7FX9/InYTDdKKGh
MIQMULT7hURo9LWfXeUngiQLg2ALM2Wofh09/0+7b4cjpNjdUEGyOkwKxTgxEKJm
T8Ci1nuy0GcQt4jRRgmYjAEYlQbmxfiP7guWRv+FnmfuLBZVxWW/WP4akGuXprR1
VhZ8eKVvWB5mVES2rCTXftmVw+CMV2y0DkyL7vATnaW9Otf6pLQJ1T0rTnNiCiTd
dWVphkje8y10lonFsiJCJeGVcLTX41RcPajig8xZe1kLIY0c5evyExMDEdtM/d2h
eGa2pN3yNtnoqU7UTzGJzAqpZ7zdyIBpOVS4JbCCXh3PwK/Yj6dwJmUmMQFgo9n1
zaDKyivPDMAxVDAkp9qjuApKsHUWcDugncS3bmmmgneFWBXVBehnl/uHEaqWJAPs
8aiIcR/3ra6qVxZX/URExGNpGnjKCoX+4N6pQy1czYLLUOWeArNCWdvZ5ha7O2h3
O5gwQAKD2EpZriDRwRQq1K1tjMK1+tQjo3HKIYluutpMdg7/tBfwgtQG+N7qP1ho
tRt+u+2l2oxaG2Ye3jEk30bdslEAdKwa9a4mD1pDH4/ioB1ebNEbaH9MPSqHCUOr
ZheypJ5ZVQ3WftjPlCP1u6qT16CC/Uv61eQzFk0IhlN+KJkTYLWnhf2SG86eBt/E
lyaY31a6VLp1Sp9+5qdwWxzqRsIgDU9kpYwc+AWyuhsVT65bfGE0Y+cztfWRF//H
WmaL274G9xYSxm2Zfj+b0mLIXUCoN2jjtCeuljP8uYTt7UM1vwG6u3v4Y0JkQO9Z
yLbuHjORmi6elO/bEEbv7Y1/8RRML7gxeGnW5xN1t4JllhsI2U0yCeNyI4dJQqOr
fiXFXkZO1USU0j6KMaNrtxmg/h2eWScuW3Sglrjy5AB7MSQ5nNzNUNVbD4Eo0RBN
uZylRiVUQs2j3kSmw2QCfn+x3vyhJA+AR0GJ5Hm91v1AA87a7kTObgyFUJPinA/9
kAfjt3o1j4V3QXOSDIM1AdANP9Wegcwwujdu5sBy813xpzb1CUUGPxhTkUzSPIF9
WDE8zOYFpjFCa7FMxqJc/HFHcM0yomDUxUe86War5Kume0K97/gTSaoG/ng/h7Ey
aKJSAt3W1+TVbL8Ht93kM3TfhXvwZ2vXN6NgKli6BUcn0XNGr4WnDDJAqThM+TLj
1wEKae3XVxbixxSlDvR26xXfwcDxfmlHtAzcFRPxHX28oi0SnLgiO+g+UEAnHGa2
Ulf4j1HbzL0BxocqMg101k2T1xu0zh+aedzrzNCluhM/SS2aCnju1hLQMgmsHQSX
sJ+ofuSQaetwXmDXTLxkFRuuflcVun4Jbg7XSWJULz499f/tdnJqTqih0/iow2+g
wewc6Sd7/6LUl/C0RHNBMVUrov7qBGchYZ46hkt1t02+3FyIVqJENiCygK71346C
T0XzpRFqb7BQOATGeMF01aHhVszBMrsQPgO6uII/OVVqMO8VL0tuK2G6HhScLO4j
OSaKrjsIbtG54wl8JU4aBiH2bRUwUOpnwDk3p6JhfFptVImKFuvAETzuzrS07OIF
2lmWOUgX20nR0OkBkzUfHoJSvnSKqiHstyK94eLWQcbm6R/QjjTEUtW5Qt+G8OHC
z/ybpOHCXcM5Du10N56xLE9p4wPgiVMBPeO5JvFQkqzmNhswWsQkUc79c6nyit9e
w2ZWaJBp91qJ2KsXSiYkxM3IvtcXRzeskjATfa3W7AV9TsHzu4OK6pYrGM4WuYww
B7yNUNh65TVufcmlXzr+pDLZd8MR7dV2GrSGGEWgTbpzb9zB+qoWTmY4bP3jiD0y
kKnNbZHV4ANFRiBIOcjadoaShmM5/m0PfYInIAPMIlrAn864VrsqhGqbqjGmawhI
7wea9itJSjZKOXQLzWQ5P4jbJaZMsXVb/F3eR+6RxBhJ0Wkq+sZw3iwJl9JJKUOC
BbuQU5bX3KZr1rnoY0l1zT65I91yhJhnZ+gnk3W66gYSw1kC6u8lcw/K0aMCMx6V
qCcY5OJu9W5wpnIuqFtbp7I3W6Gf6c3z9kyagCqABRysfMVTLaunA18lyaFwk43Q
qO5aporGLckICIyE1YaEhpcLmBt4iZfGTbXHtBm51f2WhdwCDgDZvHeWt50QChXX
bmM+NhtoMz+kCN4EcjvZFGOTCXajUSTY468d7IaUHaMbIJ+BWV4X/EIsy9PKTfYP
iIjcdS5YlwmZE7L5dyPf7G60LdL/An0oObQSjV3KAPTtpbo8ANNk++Y02QS8Lcwe
qlK3EerZeYmcVcE6IlCGHbX29WGBcKQzu+VCKRqgZjEU7i1+rVIQDqtJ8ju+7MUN
Kdo81QJVRCXRKeGwqLk1hxSwuqWFadyFcKTgSJC5rCjRKIM3764DtDT4rbAxTh4E
LvNpY9iOKvos2f+RXRCcCVlzXhpZsUepHHARtKexadNEMioxdqrUC0JUyXFeIntg
PLfc+lq0s0Q0u7arsvmERARybuuuXPhF05yICH/Y30HddPsfiatsuRhEOCWxCqDO
1ujpz2ykVcOQupwGc9xC+CCIhnbIYsTxb92BgT/rwQKNIw8xrT9SrACLoceVQRRs
D7Ai9dCbbI08q+I7KYdiC31YJHXm9OicLKEiKmQnywR32KUmpO7LxZmMua7XIMLZ
G/0Vu5DUFeOP/g0t0cHKUutbNLXl5iLPp15P0FAtMHWL4TG74tNBG4RhPTfJ5HGY
QPn8fLOYURAd0ADE/2aimGKWmesRAbyT2ObVsTDG4umeKKu1EqvI4hNtCHDmlawY
2m2Q8+uM3Y/bNeyNgL8w7fAJrjt7Umek6PBUa4DL9zblUeaKVO8mAqCz00ur6voR
9oeImB328aHkIgCLvTc99ztiFX/FivrprjxhT4CTuWF+dHbGOXUW4p0S6a9lqqHb
Nj0L0JFUsOHFoV3kUvE+Zt/Ys2of94nh7tqHBROBHEqxawaPmO9cXH3rP55ZyvNZ
tFwASiFLLUW0SE8Vrs2yc5ASxXNr0ED1MW9uy6FNBt40FFCcDgxkbQNLNa0ajPkQ
XgJBD3OMaIQ/ciQKJqu5IxgFTbq34V3H3DTun5HVtos8Thhb9Wikmn0xMjuq7WUI
TnpTxxfyV7V6Q2/GQxK1oRUXuIuJpIzHq8r1IEISqQVmDYNagMwQkpddPbvdzBoO
4kE81rtJazzrPAmn0Q+KEdEsF1VqasC7eIwClucrRB336dnXENQ3YuaMtzRDVETe
oNpUJXS7ag9hKnmF81YghtN82ufevYwt84taai93IgJze9EzyZqkb3oQfj1fDIwy
tYJbs7YbvUiYP3J2K6eluYyvDWLC+D4UuHGNHQU6WgOHzKverIjQp+Q2vsGrj9up
RkEItPo28O1e3TyUdjs/tTSIE3x1MeLUE2ftBlrcC0eMs4lHqE6JkcefLOHVM+af
HET7YmsgspgHt8thDGkHgR/e8KD3ET3xY3aGaaLJCwWnOa+bRfVjwqvhFoV8bI1e
xmJgU5Fq5rqCKi6tVSHRo0dsnTvMcNGtlh+8e30uRTgod8YDCnWLnFLq4arUC9b3
z/ocoPzZo5DZ/AtEGB+n7S3uz5acOcEEiIwW/7etSeG4Ky/KiEJHq/bsQlXxESmQ
6rH6lkw0vfVtdV+8ZhQK8rjSgJ1CenhQB3NtUD8ZbFM94idl2qmX5KFjG7btfACg
DdVmYZSnJpsMZMM5I6w4jL/pdo5v9Eh/WPxr85XU8E54eJ7pGpgCjrTTbS2b+P4W
l039GazoG9VmwZ4EfNFfej6UBX6ZE7Q0AlejjsMWpK1mLEMNqLH+29Tue/D7xqfE
TXJ+yRhg4OlecU3m6AVLm/jVZ0Yye663aowqzPW4QgSX20kugzPI0sY+QCAjvj65
f7vBpvPWuPqEOzpM6kSFs94sr6FbzUH8G1BR5sQQiEZpvbhUiVGvnS6vr7wFhCRU
aQlZ3Xcn1+XN61gHmsar3o+hGrYRrWMCdmXc8AB0T1M9u7qF+mOwpxxKVI/SEYq4
feKoizIZeSSWBw9y1sdtvbwcgCzV2QborrJ4wW7vZdp4FHk3RR45xRXOpGk7IkEF
SoihbEkf9EjhZHC/v7LQlHAVskXThEpZx/CMkQ0J3c32mWmx6iZetkQtm8CHPBeN
iIUxWrGI3GoR0rmBgZJcKH8pU/8c6iOKwlhmOOfi8iCvJl+2jakDkCOkitLY4oQR
9UX3UrUsraRb6FWijXCgO8r9ImloKpGiCaDymGT27Rd0OSxLiCWxKlPbJESWNv8O
SdK9g2iCMjXpAGxH/VnZuPcKpN0V30uyoUwynnvKsuYBiNNtgM8w3T+5cr32UEVP
aA2J4IeM90qlCnND3acaqzKNo4WjK62jhnjz/GPgPFDNflUNZ9HMEpGC3O/+SrJR
VVtY1nCjPYhdF0yG6XfMMQ2GgpyOF292Z94duPE3OFkExrVdwE9SuMzEh51cmBf3
lh8US3SD0igYTzaXMo+jsypsgB3inCyuCThq1J3hHAnngsK0XhVGzE9JwSn3AhBP
mdvV4CNLS2G6+CbzUP//PiTOKizoS8X02NIpbKbesu5FqfpiRxCRsIDM3GnqoDZ2
snvjrdxWWk7q4SR8ytjbnqRPKAjzL+sd6CEFC94tKU1KZXPMfEdn8wYrwraw+rNz
3RIEIvZZvLbWzZuVY40dNWzqXQrG+vv/LMYMlGE17mHPXlghfO4prZSjTk9n7WTW
NabTakBnhPd5B+QQoLOjKRJT0yR0j/Q2yRV+t5u3JCo6hL5SnNNyYH++3zOiYjj8
M/Lf0bWPyLPfIJme4kGMmYZ7vfrZqkljlewt2llY3FfF8HmQonwnKvZmGlSj8AxL
40859dXzb8CYNdunAgMY6TcbXLDgDCiaFGiztVHVsrpx5MkSLeQBtVccZzKgep29
jvKXAoJBQfqCAcGOq/AYyieN7rpBaGJsv4HF78iuAu0jhYw8Rf6qDDZnPtse1v9i
oFNv4rBSPDPHsuUG9ivc0lfHMbSPuSOxEoGhS9qrJxMpD0YHyEtrgPztG2u69n8M
3vjIiInoB4CPDj7i2JQcvAWZKCaMOt+AIq7bg/pa8OjhFJ3pD8+9kuDbSEFzxPrC
jDCT7MbjmZzN5967aj00/fpYqZ6fZpXF26t1fNVP6L1FIZbwIiZipgkdTVHAsmDu
uZlmkBr80KLsAB82MRYc4d/hSJwZXFKnIrzddkcfbr7nN082e4xY6NVQuix1Pmw9
QLGXP2XfyInTol8pKL3/mYU3WNYVd4IrY0D1CKmZXoWHYGtDP0vJYmbQCjF1sYq8
gYcLKtK2Ljkcr4Z0tkvr49J7WpHc6qiyuDHAsPTsVYs+so0nqasEcEUrzVIamliJ
I62wMx7M6n7Ckb956buPgX+iqRqFQkk3D8momNxvedFfCNsn2HuYgKcNVoWFAzF3
4lY1L8MVf1mjtS7FB4REtA7uWUJn+/9ucBzP00a8DBE9ZjslkQs8BbLh9ZEk+fqA
4M+1FysJOZ3XqAJp49hdn1hgR6ZlovbSAij1YtnVXdg6jOGqjoG/7C9XONBjaNvr
PCXoiFwfJ5dK8qyGmv802Cve414zfCjZ5nA7orYIVGdXAlNXrhhVRlsnHqeaEK1v
MZpX6IznIvoWQd9fORgQhq+RoM8zAeBMHj0bm3EQF2WCipYvFG6cnShstFB1KJ72
4fcyqzgrugHc8BPzbUxmbLJRX4hZ2yXPmMXrteC5C6+8Q0DQfs7F3PRf71W4Dvet
izh+4l5HNup4cHshENr1aB+hBR47Ey8W4rHBZkR9RKrD/4ydHaBqYnrjpEh/Vwif
fe9a/gwgm4bV00WWcJT2jKK97TQSXVtpfFHW9bSOJco68hnuJAjDH+AkWS8J0Xsw
ZEuenMEs2i7e2s3wN1MsEhNuJsUdf8sw8Z+5HjzSaSR2pQH4dD8bhmTATBOd2s6d
juMEjwdMzSpi3kGBloIjjg0O4tEj0Rq1goyHGtQ3OLRSZBhXkZtA++5HJOr3PlH2
QrnW5PGFBN6yyBHlZ2yTuXr3Q0AnXM7yO9PwQfwdCsOXKcytJ84inymB9Jv+DpLE
vCPtRLaP2p/S3osjvWiBYYIAA/WepchSqeq2dB6mc7Y2VWQxchvv/tmfkpOW235z
Vrr5yM3v3u1NS9szOoiVScO9khGt/hPg9j0aDRlKrtFjP2RZqlptPgzVEv5rYk6/
zFwZSjC7SKSvwpQ/SuUO7Jyr0LAhD91raplBnpKbGlRP/LSZbVv8gUsvaBmsZCGR
DN+DpKicHDG8W8kZO31483kZviGX2xEBosVgd5NIvCeX4EEK9oOfVsiOMOUvhL8F
mnIQHcYYwI1WX9NGlxFe6j0Dg3mMBTqEkq3Bgox7ChmbgZiXagqHzpamQcDB3Z4F
SsOYs/WGe1Pq0Ahrij0PWLqicNAzGgZO9BfP9MZf+JW/wXXoJSkZC/rcpiePckME
rD0IltctsKmd/43uOkDu89pixQihGvIb8ADV9Lucl9d4bD9v+QMbH8hQ6dbEQiid
Db7m61b22Qc2R2IX4CVdkp+YYTDcdKe4spbLXQKNXdfAVUYt9UQRDylthHjMArgJ
tV5/TjMce+vYq6gTg0ryoGmgjPfz7SIiBZ/6mcoSWn4jYaz0nAz9dUuppvzKDWk7
Ht6yKI2T3j9MXezl+AZRvpBeBlclBG/3csAACAfdQr2fK85Zlg4golGjefCwH9qk
j0fVZ0LYX4BSGb+S7A3ZuLVsYMii1jvuYgbVr9GJkAlkKSkmhAuuO6oKcqkDZPYm
FK07s51dFDISzVUoFoSFtgZz8emeGwMMw95LB2kBZP0ZsyjB2zZ5pmH0020rTnfs
34cjNWviEO4fIjuXOO4kF3IgkIMX5R0K60xq3AzeKAEOdKDbAc9B1En4VJSnBO7K
ahhsa/WC9pnhP04i1K/xeiaJTjStKF2+vnEl1rGUXbNTrjqt6EgOhXUYglRSDnc7
3DfgG9qeFyyqKKy8hjDNA6HJlikijwRTLwmMPfkxVlN1e+RI8Dx8MaTHNNqhkGw4
itFzn61Gs0aUuvrRSJHz/Vvqim/VtvkTTBoSNzKnvLvqHL4m+wcN9gLcT4pBQilX
97EgnA9kIDwK5k6ypKHy4eSqMBi65o8dNcmmhXo49ulQXfA3uZfGlhl01GpQYQF6
T+LunlelYv/0kWpmgj+PvZhWIhIEKVaeZ5DTf4Ruf2uGD4aXv5NwO+bxYcs6SwTQ
F9DFHHVfon9EBwp3egGbpidgiXLs+FbGW6IDuJa4pbR784OPNhCg0ZQoT2L9K22D
Cwrgoop0LC3YEVUAAYYGNsylRdj/r9US8xTlOV7IQSOMy23nYjx9oUh94Bk77Pwm
bHCktORLcuBe/j45X9XhayIRHspHg7GKspxyqnYuF46KdD2afQMv93XXaSZ6B/Td
96OexsBZVrdqxR5FrpV+zNaoaP5lun+wC/6ACDbCngIxNUuS3VjIlry+uLBntnxw
PO96Dw5qms919LqBAEn+j9iAc53YMZCrYWCIFTfq49ZZZhqrbqKoiGFuPx43TKZE
68ZSqVvWLfKqxpH6wIljJtGqFZJB6m1E1MDWN0bhtmaweQZ1wivHxr0riGMxu7QR
Eaysc60T4Yxzn2JSW9OuWQo5svUpNJIaKxkRb2/oFPBsT/W2L16mvlNYdHgYoTq4
HOkV2op7IRSN0ArwiIUky3fESi7PU+3STcjp/vaNp8VyQmXCOX7/ObclbCJ9IiD3
acre8XCJM/qVeZEJmDNa8oO50wdxNhvcq548q/7gwovECQMKrxyRzoyIz+KGuvji
yPLZ+NW2RKKaSwFIXmS261JjJPXlnI3+Nfgsvr2vUIzFE978pf+x/TiLMTm//wt4
G4AeyDsgktQ47VzTHqlnO00JbI6PNJ88zCnuUrZQ7ppQkz0aPG/XczOFOGu8bkNt
ZcjQylY54AY8PR/K3m/hsSJgp4ddYNfT0emd469DT+hbvFpGFK+if75vbluQ85sS
lUuQpNEP/+tT7jZzKOdBpXaGesA9sIxXyWw1vNUREnMqngpu1vrFz9EWvSHO73RG
k7p5h00yx2hqC+cU+47E5Jw5Hnwvb6SQYKsTKLXc4ib5ONZm22WWsxJVyn7PweKy
xTVr4/vQg8VZNwYxOyxv4Mcv6LgqOFNqLbMsXJeQ6EfOvP0j5Kq8HUnPkkUCVOBY
rhxWXlPJ88f680DRGx+5Mul68pHWXuIUWSkoSHtwMxFhE6QV3dbHFKyNIx8e+FeG
7E/51hYev4tzlC4HHySMLZ9mi/261L5XI/AT11YZ09eIoVkG9jOtHkdVRzPVJ3Aj
79JuQMli9J+DkNol9wU/vlax/zBPce71NdPSm5IFaRe7uuZX73yDyyoU12BfJvp4
gsq+XuZ4MIReY204yljC3Smbcd/tXtSM8OPEhyiFUZuxQASU+pCoqL1GeHvW1tU5
Jbw+OMkOsKub08VNyg4n3I3XXyFV1WsIaOuduKn5gw6WRUVyk8fCyXfwtg4te3bs
/pxt9PhFwuwczBVTMKYgktnNt+MJRfvMRPjLE7ljNOLUsYyNNYUhE3b92JiXaoUt
jzmwpCo/3WzH96C98MhPYUIcclogvfDl75wVqiZ8nf/JnjEj9t3l6Uv7oRQm55XU
eCuBlWOhmkjIdvmZJobkFd1BnuN+6VsaL5oGckZeiuxfybXfIQ608IQbipAIZ/yR
YXFRtoSIp/w9JJls0ZkkiHBuG+0E2FrTr2WNGtVydQ7cMY9Wp8MLSqqblpN/D+oT
ba1iJOakMIfQOi2AVwW/nKy198NN4TBZmycsrZCTXvh4ZC7j1F2sAv0Kb6W0/d8i
fbYSBwZE39hlGX5JuGALGbQtBYNOq7CHIrX7AZr6eJBJMw1gwOYgnaQMdSHKosrC
1CtP7uXc+lDbSmLzGYyEFWKfUa9Uk2LbOPap3ehMLxfdrnndDfAsTcN/Vbf9Kl5p
MPSTYBSTkew1lkUAX7vTglyUvxzPF2Qj+Giwq2cmYnr2x64NHUjf8AHRaHoiq4pe
XBRxeh/yKpHg+8JFfKwtGvB3EO4ionHHdqHmPTh7mJZ79e7u3xn6TkdXj48pOkCx
E7pIvgfY90cNElZ5bqTsohAnXOhCirm1XcbKm5Inv1U1aC1b/y1Y4o1o2O6GM6TK
yCFPxpHbr3h9TyZXEl09rPP6cdoO+mX1ngYol/xRA6aQ1LUr2q0wfL3Hbum2jq/2
BrIDHTcHmTlINdVg3tzEeNCcU8hBJs2nmhvRIjPHT1n7Rx2CnzOh8z5OBkKCYwdv
FvLfVOrTzfuHtIgmfYHh4nlMVRh6ryUZIGbvKv2X6n+Aw8RGEV+shuBePqoaGtLM
ps9fbDDuWbxfzGnsAwQa0oe9jR6vPc0LNFvgX9Fi9vDwPwI9gZsxszz44Wdg0luW
Kak2/uuWe7VT0Ltj2hirG+tw7s58zFXwb6OPo25Gu0pGm3MYi5FbAY/hSU2MQtm1
1sA8mVfAkeEOnNZvDnLp950uxvHKJKxu9qnmn6okpPW+2YZIg6rjHslYnNc2K3ov
2o8bSMMLzyhIhe3aS4Ueb/BkjnZFTmaKmkcN2+O7kHLbts3Ph9ldGZr20jJLFrwX
fp7PNBmasozG6eviAbVC//LZVlg90e00MnEqBT+9ufjzbTrK57NAcNRjKbGAQSx7
U6dMcQVOM4NifPl1r7/6TFlV1/NKD6ok1y+u8jTuuvnJbuRm6Ku+as/Ypjz0IQzG
tziehAqOozEOaryV1NCtAduCkRkHZBGXe7PgWmSIl93jqieWlCBRpWY0NHghp2+v
BUso1Iaia2O5JS4WOq6h3SnPaCg6GXXMQh4twcKYYB5E1VTNRNPBG/bWvLCejsy+
M/YTATPJ4rWdZxeVntO5e6daJQMKqQAtg3oKCdqjPQ2wP4kbYfeT1VGfBGl9kzNZ
ZZnCbiG+vls/CN3O4JkbPKrwh4xFPk9OOalX0b8OMoZGTdhKM3LTmClAr/mN4F9B
iGE8KJCQ1q7jfwVCOVVNvTOkFDad+CSeGWQu4CG0SwjaMwbnF4/mdOVl89NFRvHq
RUox91VtOGyNvWvxebD0MTzfTkW4HHpPzECYY6hWA97Q05aVJmzk6qIqbvZPb5KX
68T+HVxWjn/79EzUIAH/N0mCULKuNhBRL8jhoh2QL6s5o9JMv8G7iKpv8Mz2F6WJ
2WEThaK14oraPNfu7YfVsiBax/BxUch0Qq1VKdLLZJEWHZysWbfZBBHut6/UXZfj
fb+LokgKQ14JW8Gj57pd4irI+zFIutc6448xZDe1nbGXb7RlzwRiS+vk+TN3Aw0u
r6jx3zGzagxRFj6iHbtCGMtFd9zxM3xN/eZYrRIXT+lDcZ+5IDMcpYGkZPkg8/xP
Ob0tZafj3XwImIqTwVPSEIzpr2azqiOzO8rAdbPxsRvN/xAyCrR9k7WHHutxBBMO
8CatYQl13TknEQn57oUV39vd46TKop1IVQaMaqW2MWimtCOjZMipLTKFsUkHuozC
tcdZ20OXiE9c/5AHfVak0W3dtTNrR8tJQloIazH9k/SAcSTZmGZi0il9UdQ+N+tL
lp7BK1f2taN69Ocfh0WFQVx+cbxll1FcJtsIcXzBSO4/qtUbPio2BqEeomgDQEN1
malySfBB5udJsv0GVSADMkyQ2DIIpVNR/ScRJg0b0mfroyG6FBZF9b9jlIneZ1Dx
oupz3nqjbzqP6IbsSBph6yeQbtu1ov6+5GmgugokYJ0MGpxtHuAHpVABmst06Vp2
zjYFLdl4VXzfVWOXQQXLVvltOwxn4MnB7znOQ8Ppz1HmXptEld8uxyGtUerBZGOl
82VDC0991DxAV2IIAP7Mejdsx0YYWYEmPQj10/ehefRgCkcCEqkcJgrNbsRWiLxv
LSI7m1fdrgKRijXGLOi1GuPb+ehqWar6mW0MuXWq6IeWwRTgKEassepHOKWCSCgi
KXu6irEofzrETgHmOK8NS3lKgINwmrrjrmwW8blOP5umBkqKLqS9gHhgWxViGLW4
8CE60pUfk7j555KtpzYxRN74jg+gk+VDAXGyRLYYnaNoBAJAwR5mzipvDOre/QVA
83eEOR7R0Evpluo00Rm389UnnxlRXX3arGgBMttQWLEpK3ZdOWtgkTtGTt2vLzti
P4PEPg/gAtaRti3M86ZzkkQ3W0nf4hoNY5N5YjRUME9M+qEWij9nEYqyC+NJqqHY
3gXnFF6lPvYpx7+p00pJtk8GbuB0joIp8eIAo/J5fHrrdew5Lu1LvPfopoELQytm
kY0a7SxJC6KtWb+wb5/EUQlPCvDlffSAfxPbl8KWWrZDymzuj/se9CYNRZ30NS7l
zNQ4fvUn4ORhin53DMt+haZK97vadVlm8Ay5FgbtUgW//xQFZVISp/8qodwlBEQe
G+br5NVYqYMVZ3bMl2x/e3xvkikkp6SYzFaqT1QVd/9mN7mkgvyLNGU/23Fq2ef8
mRZ9PlJuAWRt/5QUD1vo+4rem7yzBu1+Sr0mxG1eTBuONG0vKW3NLUlMGkYr1OxN
yVx5NTzlxTQ9FRSPibXBpYmzEwGbAytd3hNOm7Xx0PcPd1imFbOrkBKYH+WCgOXd
FgUj7DMjk/MPbIk+5Bj+36e4TKOMqLAGFZL5KWpjZRn3RRW9ie4LDwlvSYmWwmq/
/vC1zQgV7bfXv4qordoxQzRfNUbTa7b55FLUSm+TKpmi5KpPCSXoYQcPnk2TRaLr
n8H3H3dLjF7iBEZmWGWOlg5qhFqnGINzsudGakAI8bHtUsLH90oGMqT8PviLrkcm
eQYv8j0JBikDyJHcF0WPPBk7yYiiIrmeK6D99wLlLQuaOgDMmjaId3gvOKXhfPcy
4ogeperArr6YTJfm3naFMAd3H5EMXANcXcdM0lsDfyG2GaUfxabRCX4pUw36zGW1
eJqFN3alyqdy6i3QMkDMSkK7Fa3Q0onkI7j5Hk5SeJpv2ARb1ORNiSFbFCBpoiqg
Am6KGw9ZBhWZec3z5SY4BhwXNmHJFN8g5Uwdo++SAvRfUfZLnWdAIkMULoXpfRt2
xpPtoz+veA4sig3iTjgjvOi8XSdXyxW1IZA2svZpbO/5fhYlBYTXAtg2iCQVPAV2
D1ksjVFdLICXPDMdwZl4Sp4cOvzITAQJzVusmvgwc/pemQ6Lb0X96nfn7RfQ9q/k
YQsTrvknAoG9v4mH8Adc0NR3DDBFcEy/0wN45EQDR0JLNyRkBl+yQQro0wUQgzo6
iTEu30Fi/Jf+WNkib0GjDeYeqPdJxvlq+0a0oblkTPl1bC/0Y8QgYQz0QX6cVX44
CbvzP2LW/nroHhAU9wRTBP25K3yZGkbWyKnE/MXdg3EQdjqoz3ZBn9bxNvrA3G3O
1ETTaei5wKXzwMCjGi1MxznuRCwCPET5bTNRfELAH+VFmflKXc0LZZ5lXdUjrXZi
2AYvbSw2i/ssn0RBgQ4Z9td9mF2fS2xMef7rG0gibslnl+r/v6n4mBtxVIOsI1p/
6/Jc6s0LGGpv5HT9MPv/NRl7RyvfGUDTJtJ1AIdyZeEAEXAiQdW4JIro+zMkn74N
QJvGZslz3ELv1QiamxiWaqRYaGiwQuDPYBO7IKi3jbO+ZORqqF0XPw+QYPZ049JT
ixugC/XXoGIQVkT4+lYiNEC0Vhzupy55wPGlNwIUMRcQ90MhOe5ikoI8b2Etwyiz
p5S0TVtL/6sOFWZS5dW4p/P1gdZ1D7Hb2uI/SndBPJhp83co8rGNs2/8CyAhpz8L
PjiMiwCd0t1L1G83gW0daFin/jOfSQenf/BQvZrl8KRjEo2gyq4FkuXiPb+7FmnM
zLd6SPYUiRRyPsJUlkMHjwNoy5V5v5GG7PpYb/dNPtg/v5GS5l/al9pC299pUrgj
71Xmxcw5xnnHDDU4XfMoDLFR9+d+TzmEd4EZaeAQ1cxNgld7Ac2/wourvh4ELuHS
3KF0fhZDbcCJ9GSu0KBW0FILvOE3pgbmTgDlB+SD1Va+jPkD86hN2jrNNPGC2/UA
fmN040iFbhnSkWntsoDljjttIjc162Z4M3NejHvL54amblkFreQhdsNKqyLtIdUf
Zlv4Yly2w5iTDj5UYB057i0Gj1wu29yx+Dh5HKeMIslzX7gNjOSDK+Zhae7SPr08
7sM3e8iokPyhHyRiY2B4Dhnl2c14cpPuxM6exMO8CDBzBgYexDzVLjoFQFqDNlFP
+x78BRkE9ZszBg0H/1o4UfA3qbRWoRoGfUmD7w6tyAOc0oDIsEn8A2VqBSe89FNC
4DFLkpKxSzjmrRezx0UvYRVPK8cPJ3nbyp+xwzS0u69VZ297hqgJcIdrEw0fX2GJ
M2YzPuH4qgcoPJslUP24IvNp35MrlyWIeW/+sn6I28hKr1kydDT1mkmSN4NEhQbl
xwxn46LVV4cWyZgl6wCy2lDldgzkhpwUIWxsLGDf3x0jeSnYBd63ZFe7Mw1uhvMp
zH7DpHzW+YXs1CZmJylMSCPUu9rjQnOP7O5JeVuJOD3rYE8Ssb7X3r3xFNQnya10
XD6nm/f8utDZnyMRQIQUlyvxwkBsKtcJ+wCKO2n9FgDAa52fN5CVIJO685INmIAO
poe0Jn9YkpKR6KQdBdUUnVJOoE7LBtTgordF8bvSeTKgfCBfsKg/54Bg1dq8tCPI
YMjC48p3xnM8Vhm9F7YAiV5WQqPZc370HrLl5fpj9t1kU88BngwGyEfBIlpUjj9V
YQ9bdmjkaxxfhAyljfRtMhSE2mz7d+ThKTecv7roATX4SSkwblBFuo9GKVXqxcaG
BiZkVCf2wtxa3XNLUI48CBPPo78DH9Kfmojl4WfBb7VfesdX+3THRn729CM9cjwq
YsslMlOlNRIVtkvWeOVIGV+IInVb6IZfBNJg2eRfkIGe3rXzSMvHayFLXEIaOnr8
Rxm47gXMh8oRtLurHWm5RZRvwB2dDMStZ8u4KXVNabc6H53v9imky9vo6VZ9MMPb
fXwgwMrhPyvv+QyblPTWZV6I8IwPyQuMBFwCKKysjFiCUkqW4rWSzECB8vSIO3jm
y9taKF6i9WSEmLzWKYHe4Ai3pY0dWcOK5AJHPKmAvvJ+i+sfSuV2jpGxkV9cOP0S
jxfSw2Uokg7AUWOW+QhNBXUE//HKph+G1PUAmQ0qGYRvVOjQdx9xcrqK3ZD4mKax
rvxJm+GFNsON4GkSeC86ufDxyhiDK5gTIkvcM4++863vp++VuR9Wz80Yp1FXm4dV
bCeHSm+V97SNJ05HpG4uFlklaotmUTzAvXQVbnc0eom4XNVvuULJGybsk2ceIyCD
8xeymiRHD2ZGkeC5prWqD9Pvo+ToGZ8j4/77uMdAxgb9L4zUtFxszsuiBSzwfmm0
ZfE08S1BFd6LgRCgDZ08TgzgoIqZwh2wW8+SyUyeQoJAKp54W4/q0vEPLcR6ReNH
CjQv1QwW4CsEM2sQg7RMMtK4y+vm1w2po7gD725ZGiUqC+p82ffHuijOlCfWUWN0
I8s+AFgOfVrGR+8QbDXIHz2UJ1E9lr0NQfVtBD7PDKpwB2K6MrKnsAjzR62GAUqe
An9ijuzig+QDvxI+/eTwp+Y6bl8vAUOFKp6lgKNoEPU/g+ZJYinod90v1/K/g4Y7
xufoRHtsPHHTCuJF6VFgsoatuj4vTm/RbbzE2gLjcLzUeaEy01Uwo5XkbB5XIks2
Gsuiz4+QMyUVAnFb2VqNwGSrqlBIdpfvrfTHPhGr2rT45KdSBdF8ZMIuqJAv0SPb
mHzBsWNhbtxP/CCjG2mSoQma8LB9O6NDV3yaTrM9O47h6Nl48nIz2qJzFV4jLxRe
rNd2EhwCNc+tcjwkzEWaPNHmADzuM+4uetAXrLBMCoeCD1Ufkw0ouDM6DEUMC272
AVx2jdlLzPCEgL9OEWeSpOLL0DoY6VE0HtD/Y9B6eMAvQp+XxMB4+eCKDnY31Mp/
EfylVrTwJFjiGPDUpuBiZCxHBmiX4SgBdbrltS5mUEvKZjJUg0hf5d0Nw2FP7WPo
IVsKa9xsh72KrGuuvuOZNX4qrbIheJwD7aMUmIzOeiAxclACFLeXkEwCVfEKZNQ6
qmfQAH/ZmFLkK4f3VUQlSXIOquk+wx6hBbqyKDRabkOcnNbXVKGxku+QSsVf7ABg
2DLujnTZq7vnauXBJwje85mxzW0XsD9BtCOI0+eSSjVGfsrl8BociDzQ9zamqmpD
PBvmj5U09lQWIy9oHiLuC/9FBK/D7ivPcO+DRiJy07V/V4CZY8s1MRgAAZv6Outk
KFz5g/2ZDESzMb+zLU06DVcMO+trEjLPiffp1wjHZMzdbb+XlOB4AMj5mC/d8y9Z
eQLb2+xtr8CwMvU+QNcDQHTj+Ii5fXNa9xHDSkK7Y0tQascEoZeSMThURwpbTr93
xO4yIJ64kBJHNX9ERa9yhkFtCQOjNXagFpBzgrjsjH3sibo6IEplCEIcf11LApgD
6LyGHrSzcZ5VHxWBeq1V2OuaPHZ+nL/HAQyvLRBPgvTb5dqKnUOgpoHVcY0pXL8u
+3joCv80APOmmRwWoZbvhUxE92izIam+MO2AAdth3sFdQwcHkdbjK5Rur3fh5RwN
Zhx5nL+zBZ5yVDlrsfh1JQ5BY16CVvG1df+8UZ8ODpo/Hq6evzvA3g475yT9fUEs
xl4WfPuXuiD4yD2NvOt3Im7Ff8ttLfUyVf89skmFGHBZo8rbAXh81gov1cqEc/SE
xZLotS0Zd+PhIJk0FQFMGqNMtw8Y0xdIWfhn5kl5PcHyjo+9DiReqamliXwGcCX3
SWUHbmqv6YUqswUQD/lldscUtZ5I5myoYhFeVsOj6G6ZMkYgfTJwu034C3BF3v82
uHKBEEQQsD52hclP6UZpsetIPjE8Giggmh7spYsyMU1kN1fsEVjj3/S+2z/0yAP7
kDIaCV9hk9HAogLBA3BcMflllHDcp/Q/0gUNYoLuxS7QDyGao/uRUj132smKIlGR
Z8EzUUv7Ra9VOmAjs2jNOaUg069hHRqDje1rlzR9dwLCVruj2S44mIUi3JIUG5EO
zJe8A1KfpDI2g3sQL7xufFhW/2WoNawRFD+vmLVkhZpIWjojCNcwbaN18YF6sYC3
GVf14tnWs56XrB92cRLGn1hUDrYhTQAzQHjM1Gfw5SZqTJVjvmNpsnxGE+VQCKWG
rhZVUbL+juNFX4rDTldgJJqxVollkOCA+gDo08bNbMm6mg/YvhCubjMPHWQeHRym
P88fIoRKhblQpoPufjGE4ucq8vyM6pBFV5fZFdb1MOpweMvSxcisAXX2d8Zvd8jT
3YBA33GwjRYIdNSsXX8KLdjyz5/zxCxY4BxneRRZ0eZCgrdcrFcyjPUzrwVd8cGl
1t2kfHRfm1pNBRBKvTrv+T55EPdca3jfKMogiasuNE8n6bHF+IqiDDmjYXm1plpU
wMhAyrQFAdMh7jhbwvquWTrS5YRPu3vsqz1RqnG6NtxQY+77N7cEvC3PyuyOZVU9
Rl2pwBZANH+u7PW7vTrueMk9tQiUU5lnIFFs5g0I8DxwTcR7ExIX1r30W4H0dpuA
fq2i5Toqgajt/0SWYCzIzi0ME10ZyXYDyaOm055UWIY/yjz5Ba6QgYWcUhl/mswr
8ts8hBRxzWICi4cTKWJNH5nh4fE/8/cw1SPafpbVUAP0BTPvTiPJAek/IcX2F4bm
yJPN8uY0dqp/ml56fjO2dHIPshv3Ggn3UE83lylCQ9i4N3Z+o9IbuinlwpqoLQmZ
KO7Rm49UANB/N6tSJOErivleNXfo/9TMdkr0X5gvzLEt+2+2mOMeEd4J9awpRz0o
0t9PwAd7zF3OB++n6NIbLMzn/iECnuPuXvFJG9SrLz6Bg3o8EXVogshJ/1PghWh5
A/wg3CSZo9iWuy9mxS3+Z/Z3tXrYJzp7N59jz0nvJnvLritzy29xWs4LKMW0Sffh
rlxw8rEQH58IqEsXm0zEh2PMllOLSS3Q3d/K9uHPuRtJAMQHQW+a0HWeFB8xyhPu
TySA5fC5OZRt05VB5Hl5q5sIw0dJNQN2c4ZWHus1bki1a8JdOo5/hAuIAicjUPQF
zrJHuiMINkCcbx6tbsFNZi9CuFnAQs1ftCJGA9DRlOgwfnU4M/suZJpD47kA6po7
BuHdFyQ5hVqIiEPXlwnhL70TN2GXFGKmPkhT8zcS38WTXD28lfSWbTRyoI+Jh16H
7EkcAsRgQhAgl2IYx/hsZgJItVvh6ZsNufUX8ALMUHNaGzhO/O4s2ev2AyQ2OCdI
wbXFCuu+BdvDswZaPUMbcS5JTgkpk3Z0TfAItb6r+Hj2cnP1EwyLYOvzXJPBLTcQ
5q2bDrXik8bAV6v2naVUPFjH13OpPDWyeZKbW/GafqOJOqF1RtLKUcUkRcd0ivvn
FRsg7dPAbGb2WVa60qlz5Axt/P24/ZdZzekuMygxryrLXotorcY4dwI4SI51vJgz
FuPAl70+/FnKg9u2EW75PshDGtewcoWKdXvGEVkRWdcuum4GhaBt8tG+1632Rc0c
Rwg1HdtgCZzRsTBNdX8r0SEB1gIra4extHzE3ioWL3c7xEsuuwRAYDHfuJQBKz9h
ZUN6rW3Wu6WijUKjq22RPHKfvPXbGAs4xTX6DEjWTuOApmudf2wj28YgLZwGEGfc
3pmc3ncfqJDnLTVf922dj2ASazgFi8bAd3S6cXjeIVgwVRLj6Rlg/qIjEWgKys4l
heUae6K4KGW9vJLfVJegD3d30WtYp2x2inTurw/KF6lLDiVHK7cECWU09rzZi5SS
4P8A1UmPiUUa9KgvZmBZ4wUokSsM/sbokZwIakaWb4RdJvuDAbI9fC15sa/WhX8M
72UWkvLu6NpO8m5uuom7XN4H2pPlBmPbQZpT2Yltn3/cfTfoodKQ1BD2vkGhYg/K
n9/+naVdB5yEiT2NVFb8bZ2dw9Guq9FeuqyvslYtn9wQndDDrzr5wSJ/uw4WsoMY
DQhphh7fg6zzWMu12XcNotcJ3Mdu0H7a9OyBabbqEmRcZ9KsFGolz303wiNToU3M
2TVnUQVg/Dx/uVCXjHgAuiVp+e4Zwjnl/DaBdZdunXGY0Am1s2cg3YPBXSaY1qLT
eMOuKVkaPL0raeNJGT8fWsNNraitMwNWUd43/5boLw24iAlB8xUb4P2ODaL6jEb1
saAPzvjSyJZqkch8pMFISsPIWYpHm9N45/auFoP6mFxH54zN9awvQtbJO5pwjdSB
zrlN2j9YpPtkUBOECri433ZVGpmlFXK69eQqmY3Cyjlu78pkZ84lU/UXkR73bD0c
CUPIK4jZvk5mjlIoFmpemDeEz3HKnhthPNY3SgOd4pJCbp2Qnr1LUu78EeK0Apla
Yrkih/FNqav9xoPllSOLXNWVkXZWJUZ4a30DSPlJeBKz3OE6/PMp2Ng3+9TipedR
pSLK1lEarf5FWNky08qcNjPEp5MZ/UH3pL1M2xYCdxlCaClF7+7hmMtYVqGfDS76
+VFjZSaSOOtADQRYSLGlbl6y/gQAxvw3Jw32vWQQYGYnTDQT0Q267Rx24gad7i4A
2yaKDzf8BiHPo618IaIOwOfKTbXbKTkb15lDSW94QB+9JRuEMHolI4eemPX5Qf+p
iKa8gB5WoeH2N/FMjmBJzz40OsKqS5XYwLKf0FdITVNimpZhXj8Vv7KYsWbsFJTX
mBDWi2YiFvDVhMktdOWhj4XFGE/N7VGpBTCcbkJSnhtHZvkz6gV6XA2QW8pMlIQW
BBsaAjcltkOmmFbs5b/D9kbzuMonbUgWjPWJ3eG5ncyaaEBe4GAIQNs4ohB6wiXq
nM9eIfS63710Kbm5IplYd2jy3ayWeg7yDmVMXP99NKfNwnGJIRaaSu9XpeLLNTF6
xAFdb3NeqGWU0GE6Yw3924OGqte3NT+dgn7xUfN7o5FKdKSuW1FcwsbMse1uwSo1
NIwx62IaKgiajlgiREZPoeDMTRbr+O9u5QW7T8kWYIQaHQRwumPa+qrHD8B5muYL
2cp1COanlf32gjxRpdYp4Su6eG9Pi382jV5JWr0UUs/NvJvWxVmDt6QMXzBEmAS2
OYXjjy0OW2szBwf3fVy4tGotzF39A/GAyWA6qYSptJtF9ihG8IvsaSvdTb7UWQNs
yxvFVEBoxmUJy/Y2uTyCk3x+Lu4roSTlQZiKkZHwCXVHhCgnVOpqGp1UoG25NmkX
KzruLtt5UlLnfxpgsDME/ecUYzx3+ilhOqmIQAK0BlLLS03CYBK0DDYGEA2o+4PL
1s6BGxh9zoNJPXQEljq1HkfxMY8lAjeRbKPkJCvXgdC/JfujBooeiPGt7q/5xL7r
gUZZunoDQ2pInA7BA8U5mOMkmxfZAZ9kKFM4MCK75mfy3W3pWqocI++i3hR0GFS6
LSDViFghJA9yH4QdSrFW9QPJNZINLeJdtTYBiWrkMMqiXIP0BalVre05A+rqj2mI
mzY/IdPlj4aev7j0D7l4ESq4+xxJ6kHDMuTMM4eDnUnIyZ8nOt8UzHwjVmC7+dL0
dTxsFdLV7JoV3L3Sz2zIsMdD0UU1zQQWVlOilFrqmkzHiuuWwbWhW7/k8Crfm13p
vIrGitYpybjFDnHKx+Gz4AqlTrxBiANj0pl0AU0lfUjHYJEhSifq3Try4u2m4gm8
n0mPuZP6NcQ0TYUrEkOaTVgXyxQWz01DgMZ14SxC80aEy642kip1G1VxImraAIj3
kDYs7fvTmhEnBoeqEAk00n0JpltC+3fqXrFmimwVpcxiQ/zLPLzHD4nTtH3ONHHf
29sOpoKkLZNQooQjyEyGmtWfEa72v4prdteMmyDmvIHR/BkWTQZRi93NqFPy/8Qa
O6EBHmu1i/AKRaQeuwZ8o0Qv+WgrhGw6ROghIVr2V13m7zOK51+5Qh60ahvu24xP
GPiLc/+wiExzH5FCoelC8XkDKawn4Z3J/03Po295GNJTQOKyQkcn52fecNO6nlV+
B1LpaOl8PAuzQgE7EXP8kworiE7n13zvsf3faQYIjnUbJZAMfl5cw1CWrcTG7JQc
/FkET/Oe3v7LKlJk73s9CNTb1Ylqo4piL7Q6CvHbWtIx7LLf3RW5suiuLKBM/HSs
XJu/w/evByPfomCHK/oKYJOZuohdJrrc21pNwavmoCNe7t+aH0vBoBTQtNgOrQAV
edzFQFfnV0fTMUoXe9n/1ljncMPpy6giZjrUrOsAdnE6yKycSpvyrKDP2ue4hor3
NSZTWueMRYAOcVjusiCeQCcxDOksa3wK84cfn05NIug7X8nLJ7Fkcfq0qc3/65Oz
OC9IWwnY5X+ONVScVdFFIfpZ7lN58lQ7noyYxrB65f/phBkAq5GOu7tBKyuBxW9a
sdW9Sf2EX6xg4U7EletONMYJgjldJs4BKDjDUhXFLb6BlnZJvghRPh+G3Kip6Oo7
KGjM5E8tUNP7CVZtYhsRAiIgoGYJ8jNLQM1v5XTy6UkqZL92/lSMIoNxnBlOAUzw
KOYTZMfb/WZQM5FPAKMPdGVQihBJTqaXYc8mB0vbndEPBTc7yBDlzi7t9eLnf9GP
8YR/JzWkPVZpSIMD8Pi+shBm7uCftKMBmQArjoZsZgAHonFomVD3GmiDt660MW/i
JyAznvAkclUzzsmlz0a84DeQ0ylqDRVQni/NcGN6AXJ5e5teudJt0WXWnp8pBBpS
vsVa3RyqRK8ixMIWzowAt6yzrIhHHvVeKMvvg6pj033FFY2Z6EAQ62uaV/9bq+pP
bxFQTSyrg2tw31qmfdaSfdzJlb49rAKNlfAHKeq0yN7XA6Opy0AbfQwJuQMCYqPb
77ziZRwHCD+9jfkDNrKXzWOgsydAAAdsOK3Mts46CvadkX0UQ8xvwwlLTqXrj9CL
PNPYqOHGbVlmLcErj6QVcFr1OLqZedOgCe0hjlBNY9oja21kqzF8NJWXrCkWbIWM
7a0lAaROKJmYl73wNhR/0yNIbWsu2EDfTb6wWBqOE5sRy4S5T+SY8BuqmWCAUFPO
o4GnJndyTaOTI7xYZ3Hvf8dja9QMkJjHk/uNvCQ20app82qUwalKCVONdzDWgTm6
lRfuYFKe0uZ6ZE93EEJeYZqtdUtBXbx1P0HccAGm2KXnYHDvDbX6TLJrSicWRixE
zQBEtVfEurZwj4EyJlNj9Dnal/9v5OPpJkatlHo+AwY4whIrj1FZO73ZhX2eFCJU
MKY02b0bdMvvnzangig14K9gL8iTdYeGz3vFN9M6olwr1wxBzK6V8IFYcN8RM8FM
AORH9Z+sslhJMDXoK1xulTvFa1SlqO5t4AArELYG0qpXRXGzOVm8MN7DvElUh2kr
1t8wEB27oNI3BOjDeXx4uD+WpqL+iimdGbXWSJ5siuw32vhD1M4/LcDLA2bZ+AEE
SlJp00l5oKer/H8KYvMo7jz5UZc0WzRrzJXmF5uPs9jijQEcATat+K22vwRs1y1f
ZpJp3e1lhsJ4NZeOKVgE+aDK71tH6Udo0ExvBEi01ByioKGUvpnLalKXrVavKHtk
/hpzP+Ht+keahKX+fQ8QlmXPEfaPaNuXcGvcHHUFqWp7DfSMAmPDJYyKEFh073s6
6tMGSb2XeFgNmsdiyS5SK1iQEcY3Gg8UwcO9flGqNBUTyqG0JHrofbytFSwMqPxj
SBCap2wfaWnLOSAStdbSmzyCbL8MjIiKEpI+l9IfZpqBGYexGMYM6jB4KnFRDTGW
g8SbM4G5ssFjN9suUbV1A3EeIh28X5LEdQDlvgPItrUjOV+y9kJvBTKUbQp2ujb9
8/uJgoIxCRI8pKS9uhOUdgbzbkJSWpk/qPFM/RQRHj/mZUsAgRaxqgj9lreKIBTc
GW7u2GoxjRv7Bh7lSbOoSdsMKdj4SRTNFM4PchGFT1JWp+sAPwKGezZ5FiPgmYRk
yhDtUkLaOKn5c1u9RwsfYcvWacl7vsiJRAawm0cEjUSJyFHEyD9r613FuSXHaJtW
4fqtwxdEnNeLBn+0JJ+0D61r119w1GMgEDS7pLx2fnIuZlIqExeEENj+0DGAzBMd
vSdt289dkTzHl6CKdnFkVbxkUdKaTHl4aNUusEsQ5Hq0BcT/XALjLE0GtPQnUDya
O/bvCfal9Ew/rsb7vgh9Uqe4gGW3yFN+C/MeSAgwhHKDd/y36Zzn4zljoS8522yX
v0u/gLHmooBi8JzmXtbKRewbU0sMJqk68F63wJB/CpgSBmlRbCzSWBiC0sdsXoBM
RS5gmix+dnki0FITwBZ3xCB5ZBBIlHDgWZRnIO+4hH+4M/dNkdUfuUjVjwSw7Tv0
alUfoVttBXUgkKPnKTIlNYG5zmndEXddWC5Vwf4FXvXmMNRy3MiLhlyNnzuQHdWs
gZmPbOTX863nCkrrKPlt5Taq40fteZoDdcwdjiqfB8y3Xunjf5lOhLyVE5Bvxw3q
+tsecmWZUuZ0KGvsdt1rJ8SbR/aZo2vOvYNEST5sUhraRX00m43J0lU1gs+xDs83
UDPbuAqNIB1pfXoTYXWeqbQ693uhalZcBEvtMJjAt2ByomlsAIOVD7Px1fCFH+dg
zjJqt2sYCa/JNH+life5XN6KN0ofcubo3zCl4yNmtvFNwiE1Nq/wPVS2ltnFLwS9
mYBs/dDoC/NqT06msqjjeAN2dpPlBn6McrY3xqBmhZzkTPSE5AgUdMi/2LoUv7Wo
v1xA0tn7tcNXXpXGP2B80UTW46vl+tkqRAMsQ64cUvEEna6towBoiLgTwe4bwSzx
7bDx/5yWNOK3n+B2u/n8AlTHPIOkSNJISabLl9wZIZE8wj9xWsos66wqTYAx8P3j
bjLR1qwm+QgDk997ZrwBkvn/NwwDM+vjjBSheAacCH2rIxThsTKGJE5Iey1RLTaJ
8I0GSOZkIaOP8HIEEcQOZlQAPHicYkS8yXW5KsZFOSfKgqRmgEm2C2kmbwF8JLMQ
q05K5YNx/gOulT3lPhKi94kkYA+gLB4dsh5Z+wQl5RCPe5eVaDcsthKukoi1DaqA
O7iB+RkEvx0xIwzprRsTy/2exgyrQ9FD3uo3cajIbCdyKfx7EaDRU37zrVhKnkHT
4qtUK1ZpoNTxe8urPuTTqplcgQrs7raFwB2Nhl+cKZVlevEvbCjjeaS/OfnWVAw/
UCrJS7wE1EGgU2S5AruqirHj1IXC8BLkUmy4TZJVI3ySoKHDlZLg8CYO3/n5bJOV
dW3yaTv9Q3VhfOgBY1YHYsRAe3p8BeBJ14uKWlksQe4ah9p8iCCjG08NQhJMktMv
PpEdklgFWF6TammGNjxM34hUMwft6nszF0vVy4g7XuUDbEMxpY9qfYrxBOImVo+8
CgyHaI4o96lOqgzoOJNV6l/13dMSfzIiVbmxkY/RCWZxwQkad7kYuE4mMenuTVoE
ZZQWAojaTfQO7PoyGx/ubuVsIgDKBApl/ebsk4CG7/unm12x7/jYcKkU2vszQEvk
/Dn8NvSYZSD69IWUl1is2TatkZuWkwbvlZCogeuudWAqQg3jeb829D30RsqVT/fe
0NbrDqTzzqid4cFjcx+ox9F6fdIteMLFY8bXcwS+QBrAQLonOzDLx5qzBSIW0YuT
70qkbVlGyTV/nx5OrDp/zHbzo1avF9jIumP9lABiZ39ZReDq4dB4NXagZdJagbpZ
wnEWAIx9adTHVbDu218puiW9YqRyNme9ZO/oqwwMks8CnFoXENF7OlQPiGbBXPuV
C63jnWnrhbyxrQIXacLa8eZyyx4r/U5dsT0GloO2tbWbgewpqZpg2Z2CfR36HD3m
C91RuiDk5PzrW/W7MP/Yu2m6go61ASKiGB8+pMhXoH3UaKjMVMuYaKZV6Jnzrvgd
LDgxr6fnjkiMWNJvtW/su1x4Il47hcS8XYTD/FUZudpB6fLMYAsBc4AWdyeIUrHB
iFz+qsEUcA64NTUEIFa8X92RNHEx/66tt7aMSnzup/nmpJ+zmmpZsrVXACds+suU
3/eHRFk/xF0i/7IFk2csxCsAWk0+t1IHgysDxuvTYWGuFWn88Ggy1XDIJfHiYVnj
38fNTSQLIqeDbYbBSt1hqBqnO7/mDDEKu4bXxI0slsUP+X7CxZCRIqZ41zqjUAI0
8p3BVRLr+v+08qiOlxnWVpcWIE1J2smHOLBX+//O30VHhVkBLlofOsphS1rH5Mtp
IisztJNGBROSyeOsLepk3s1uFXbyNm7ylfykA+zaZDDX9wptbhSxMlhN1bbGNC2R
Q3ZJ25L/Ad3Zp7fEqlUFmrwPMlKYSXar4gINYI9SyHiaVM5qk855y1KARa448v1Y
C2q6oRasy3+N1VyBZ5T1VUhNsnPzfgBGYgU9TP6hYKFAfVyUjDHl2DDn5EnvlorJ
BDZg03imUFkdSp9vgrEUfmmWncGN1I2Rli/CFyi8kebuBkHCDRvPW5gNqNKvG0zX
DOawoOMRS6Obrk/CVLPdxnVB0XUbanQK1Rah8tudbZ1Rv3FAOwQzNYSV4b5AzHNf
q6wak7HS3f3lNFxLTRdw+hZn4GV1A/y2foDlKrhoXBZ+rHxBWYULfe0jYWZc37Qp
VDJz2K/PwNwZJo0Zt+a4iwxX5W8q/SWyvvZaJFnmxKGRoN3KSvV986K4UpNaKf6g
e84GeJVNKBHXZS3oCdaFGRpoJYMIklSTWk8XKOQOL8se+O5JK7/Xftldyioc+tmo
ZB/AsiqWpxRXb7Cd4CHDzQ8dT4nLn8XHJCsf80RZPH/uce5dahPO8sH6ie5ykkh5
ujpBnL2Y2J9eE6Xi5CTooOtJpnIsTZgwnh0e2esOEe1O5d1JzsS9KB5Yj0FOt8uE
UgGgbBD2DdnnvrDerOkAKBCtZyFviVwDIFXUTaVYYSjBVmWG0Ln4F8A8cDvnCSu3
BDCzQayPx2VpGRggJPdqUJTLUNUO6S41b86IKtQ1nfnj7uuL5yGOxb0OFPedhSPK
2RAHu2bC3VkMfz6dv7t+LY1siSdfBMEi8pcSjqWwoTrpVU1uUHKX6l+dco2ckimb
J4ApSE9ZQ+YyXvxxK9japi7y60I1073Vu2pBhgSNuocC7uuJ3hRq4Xljg5wULh9H
O41L/WKjzqIBVN9j/jtrzmC9tSK+QudcNueue+YPhM58+JW2Io4n74jSQ7iJ3l/5
+/GcQhyzM6HBwni5N+ORvtHvUgBZrTNNt25edngURGDjt4mXncX3USUrbf5iQBNP
0lzHwniQrgZgNy4NUBfoQiIRcso1sWwTAEMTJDrPC61Zs9LuL0ePH0LZm2LUJaSs
KQMkfjMMamXyY7SK2KyBCHybXTr95cWbuLAs3Y/g4HBN7/EWA2tHaFE4n4qo7eYA
3iPrykRu+kpoEu/iKe3pFf7YV/4m5t9nduk6rCJx6mEZifRNOAm+ZEzudmGQzPc7
glPdi+Hj1n7fPTIhO1sK4+OmoYXOCstyBL53VCEPs7dn86z0OzehjxE/IUe07pS6
7L81DsR4RueR4QWoLPI7uRV/0jS7wbZOjV6NR2fEzMmU/+8SxOh9DEpPF/cIRnIA
MfykfvU0bK2N+HWPPGUMpm1cBbS5R1m7+3kiwwPKKfrQgKaq6aPs/RytW4hC2awe
t3/G1DCNzvmoRKGAYa1KPTlPwqr88cYz6rSvDKkieF8o6WH9j8PZWXWW8bYHDu8C
AWAoL7zXajn7mDxFZPO6d5e8jeucfLsbl1/OieQ9fFMAYnWuPFmKV53ky14TKCOj
numLrhGs3tgZR61eliodL7DpaSr7j8OybbuF+sx265nN6BVWPap2oNQ5R2I79B0j
n/GvfuxxkwvBlAG60JBJTwtYrekbOdArepcpfunuYaaOsuNkC7JUT4Hc53Qp3WBI
0KskgrutKDBbTau1a90EoJMLAJ01qd7vi8WCUWDsQ2yfnnEu75KlAj1OMPfdx8yg
pHuagXRBw5APaVjiYUS4Uo8kDUEaSCDLebojhjGaCNmeiGZ9MpZHp9O3wxRpTYA6
BFbnxU2N2lHmd0RGquWpqlg1U0qz9WittOKrQIyefH84pXnat6K0RUdcP7tk1+fb
3kyuM9EgAo5LRdx3rBP4ORsIVcj2YxT5fNtSKekOGnEKJj7G1qk1gGqWYOLqioAB
jw5BmTqzOLwXUrQ9k5L3SROhkzK9WqHdjkXatW56EH069d7q1uKzutbhMZok4u8E
F7RhCT67aAaHo6m6nBedoLi849LAK/Dy+mKNqsSXW8iCA13a6CCwAvT1ZCZTwlSz
v7lsL4f0zCCnj3Z4Rb0peKqE2f4g3M674d7884AadDtaMTFVHv1AnlG8R0jY68qk
Vth4htPNjqLGz+ffrc13bTBxyk+rvSosUn6Ck2p+0pocTXaKHlMcBT41fIyl07lg
v6rAW5WBn6Fvjl3/Xv7f2cPkzyMyrWg8nRr6jtaKRHnlcXqbDwhzIqCnChqCvys5
cZh5XAdQee6KGurzIWZp/41o6KBbMcTIE4PeRBvRC8ntZcGMUp3vXfebjp3XN3Bm
MKtdb313vgAlhv8phHAke5iFDjmBPoZobdCF0ospQUVIgH9jKmzEA4Yky2yFl0zn
6dFFo8vbHZNgV+0YieF53NRsgvjeV3YWzjcUiC5j0c6G4qRuKQaJamZAdKWa/+XY
AW04hwIPFIc9uE660aeQsX7vTb7ZquGqhGvT1/SllI36R4TLZHBICevhrcA4rWSn
T0UzWwDyugV1C9TzhNNInOaoZIBxhFoNjAzHxJA3JVVaXarxKlAC1FGdKe3BkS47
bhVyh2RKaq7XIjkqMXqXUTYc5NuihsbRHq4HzL8ddI67JWnYww8Rb0o5vMJ47epS
br1EYysza3zXCKpQje1Wg9rWp+Bko5z+a5I9NRd6xPt67Jp4GQOuDkhEfb1pVzTo
Hi4MojzmBuFlLE6hbjvMJIFUEoxNJDKCBqP5X8mzpEveqYMeKHKLxUD4oJTvhdPu
1jW0WG01Xr52t6j4dDgIzGOn71JtRNDZo7wGgbW9SFJqNNg5/3N4dCwDzJ8FNTPX
w2+IXKOfyfRd5YSqN6Ne+02gkrW9cG6Yl0lwdmDGxXLULoh3RCwAaQVZLjW5E7dF
vBisE/oCcCY/uW0K9IBZ5XOGSMqc5wqpxYkqsk0rHJol7dsnaE59zzDbi346GHOl
jvea0qF+yQ+JpwOGmtHzffYmxzSXtT/647UiFk0Yauu0oeaOCqpAapGDUHCAHznl
OexzLnPE90QvQdwaDS4okV9W8tFPgqXyovFIDkZ+JJWHdxdoeQfia2fowbA7Oa9t
VJnqy77qXVNaPsdROskiEi737dkWNSmpbY+Ka5gq8hMjJcccjItsBFTc58ddW5jn
2hKEgKMhB0wDon0/qBgGLqDqGlBWiqtv95apdlJERKxa8bfvotwslxKWEhKf1PMh
8sCpirCLhcz5/g5Ss/QyNrSFlFKFKsZ4tHTnctbz9eiFZuuSRv/BZ9z2v9UFt6Vd
aWIJuJqF6sWMdov+sIIFio4w/g9c6+2XS/KOBG6/PSm/FXYlNFZLIklYXAUk8ZMd
jDsPfKf7nxone4dRI1du7KAFftE6qIdmeF0+qIIaVtz9Z7XxtlEBjoEUcgzvcWMN
WevbeXG077I4LT2TjigddJtSlazO+UIOO5aspFBRf3qdwZy4ABjYpgN6goOu4WXq
oOmO5L7iFXiNe29KZ0ma/hZabgEBw9bnqatuocI/Xad1KU1VzUuVcXBWXOKSHzbe
LPz98zPZAB8KrwGGU7FpA4jEYUSxpHuKOjiCNIKMnQDjhDDAL8yuuckfnog184j+
tKF228F8pYi6DGPsXRZCVcbBVQvOQIPKGkKldsVkYKXm5Gelt6yyiv2tP+ptvdUT
5PtV+wtysNt2oDQe2G/njhm9Dv/L5+yhrGq9Vw5FgO2DQ34QJoiUTFY7w5ipD1+P
SJHz0AC7J00vKe+9HD9iMa4QyKIKLz5FbYOzdCMZVkTCEZBNQsLxs80QDNtUemTK
W7yQpgG3uE449Nf82sclS9CBQ8vV2ogu6V26OEkPkRfTO287AwYDOsVoyJqK12qE
EjBKibwyMWAjorQFXcOt6ePIwNvILiLcI11EF8ffyewm/kcUyKHVd82T5lCN5yNI
Lt5oN13u48od51S/x87LTDwjLmRG/s0s7nr14Cob0dPhaP+njj5X97qKfWq55UIZ
CkYI/OH6kli4lC+90jAxLPDGs92d9IMKl0zVYrANBrWcKh0UXfkJsd7H5M6CAfNq
wSdLDjKON/pn0q9EkNYlq5T3NV6ApzZdeBDrq0vFwWZPc6IgLjGpt6KuaX9L/Tbx
JBEYGMxmrj/zHRq8xrv8EzDvKeL1JO3HP8MCr3TgGt4WClNqole5go/O2/pIkLpe
/y+hCTAxAGBQSO82I3E4fbc7gwldbC3QCB2nE88+xWfE8yqx+mpKUXbJrYMZJWOI
SybQ++NuSYRkvN+j8oDEzpAZQgpbRmTUMkmN7ELFZwjBWHVgni2V/hKePDbeBi6Q
i45oDIAZDtyIWq/oDhHp2NcHeKxWjJ5wnbCPVRUbWmH9778t24SoszfdUweodZj1
0xqRBzisPzfKyLvXkoDlriN62AXr/NNxTORaUdh4cR5rV5W4lQAI51p0MCUPJMaz
b9JNDShvu5Q1QXgiWMyqiW4D1R24QfvjZ4031gfAyIPwDOKOpuDjwtY2O44/D9FA
bZOacdW9950I4tr+l8itpIAWRHSmCrR+dR0NUbkjR1kPaEDItAmgRrgjL1CLBF8F
PAfVr+Tn22xqVV1YtRiF3E1rtRSxJ1votfEbg6itQ1Hf8R1I1HyqCTIK/wfLvDxO
B4E3PCF55d3F8DrJ75RWdmlPK+tZCNijPHZc3MeZDIyoiH2RLruVqnsICzXgJYIb
R52BwnWr86nGCxI5Yuo2bLysGXllmMZvVerDJ8tEd6Cocq2gZIpueoHxOpzRcvv7
BQAFuoaqVqDZWM+HzbadX8irs/NsZZtgeU+0wZXbNfdAFOSUxXwyrslDNwp3+K9k
cC9vwM4XU3Gxl0i/etYZvkJN4Nlba0I2kK4CO1UfQPEAkB/hPZDZXwOY5SH/IDad
vwz2glmGMXl2OEV62bHR+r5vUWiLHKsWe/b8UYWfjEOsSuoIYo43d/9zgJ5umY9z
D00lo0BjsPy9kZrCX+WR6SQfVlB11VXw0Jn/xGIEYXJNow8e3tvWhA6gWK3eOteD
3UmiyqB21XdwtPNHfpVAxCOeICEfrrim/VUpQVT9xKlzeuA6NuT7dr79po+y0q1J
ke6PYWj2jiwr954nIu+5UIsMdbrAr97+woZTaGrPurzu4Hi4w/xsQLSWCmQe3g8e
yD8tjGT11l3K/swEvI8pNNf9Wt6WsGOo+KPgL97dqZmhDntqJxa2TAT6SNO788xx
rqzjUlz9evGWEtpsmQQe5WUOhNwzZ63uJS71L1YT7alEhSt73aVnlQqLqxW7ZS52
bIKbnCU/siAIvaXh/qhDUsfrqTuq91t5vTkDHrhYZIZ5XbYvZWDiKihQKFiXKbpO
VXunwaY/7vp1l2MLrGZd4Zo7i4QlaYJN6ZZfVIi9/7cWZkYY38Ge6p0XicDjHU+T
xwoRjv/PZ2Yq3+lstOxEte1ljQaZZmaiiRXyRSgjct3yvFP0ZU6YaQ1ZaV0Rjibu
VAkwzxSk9KdaJak+eRtds04ZpzvEE5cgvtNTTEZJliaLQKVA5L40tJ2eC0slv7VH
3gaHK15RyZ89681pdIiE+pPzdGYgnObYc2Um0n2crONnCu30kn6vsKD/rr6XE4H5
PmjfV9ii9AO8WHm696b1JxQ1wcrA4rbx8fQoFCYE2ndq93W8AEihdhYMyTgDpz9v
XSxj7zqrQTa5Q4w/f/7HrvmPgYpKtw2Jx369ZtDuW1RYLDBvMCTyA31Wp/QDu2rf
9HcHC9KOtPLB1tpWGFF3gADS0NMLQmB0yPpOubdr5oFVrDMxkJJx+vChVQvjoXN5
VGyunA2Qse0YKnLp12dYkvkEm3AZgHXNv9UO4jiXJm0F8m4kh0czF0Bcf4MXohQs
2ZcuoRpcZLYfgqpTZKLQfFkU+CXNsI1UBjfGTry0oDSNRhH0Mz1GspsdE34ocxIH
l4561kfb051Q0Gjb/S4hYKNQRitSX1xreVyY6yF56ah4goz7BdGVR+VjWuSD1y8u
1Vb/zYlHScoKJao7hDIX9/hErbK6orx8MkgG9vF5YEMCOr8EvB/2H38ZWXbZCUXV
uD+qtZnzQrtzmkZ0MP53y4AUSub+FZHZf0MoEOLKnvJHGDgVedlk6HkkulZmjQ4e
YxyxrWR6V7f5ut1z8uBrL2PNaUdrhy6P636BL3PW+z302aBNQRWulN8kkIRXvydL
hFw0t3nz7RZWRAhrZjULy7nsi8V20dAWdlontEIKdNe0zzrS7FdaxgC8B+/XJZj3
Y3Gqrq/ZzfZ+yfV9QT5JXX3OE3pn49BYtkBBxLLYqowR0H0WKIQlnl5DEptEtP4V
w7J7EKDs3wSaQQrw8fhFrGxoV/Y7PPJ5j1o0XEf6YSZlhxoZUHNooWXUJQCNv/l4
/poPuEjKTPEwLteJixEPh/VNK1yEkeQtlsJctQhV39B6XQ5Khb0YZ1hwl0tjYX/M
BuyqAcMzDCzjsFmBRw/PpWbT32Nvuk9WAPGBSooIMbbvrIgFBA7UfYPcNIBxbXpx
4S6OE5tl8R6ju/ALL1jta1XsZbhdhrlSMkN1KzbAKyA8wPczK+rroDjOkvDk9fUe
0agfabZujr+QZYDrzoFduygCderV3VtQ6Ec+wa+8sRYTos0cnWq5EgWo6j/q7RPb
SKv5pQcmUMEFik1AZG4d9SPMex/Wmzdzw9QknHgdqn0aUQhSQIz/SW2yoNVZKmah
hIv+/4xq3W0Agkix3ITb2djjdEY3K4hCDoYlIBU7MpNnBfF+eJjshIq3hEOWzp5q
Fp2k+Wi98hNF2ZiaFJwOyxO2L+lvjh7hO5+LS/C81DhnjZZWaKVn+PUrDBcX/IcV
tcCVGt77w2pOc5mfVhUF46tntYNWhT+SCYejroyBWbiQwtyg7wi+1d8kZAfozUMW
HR1w9v/wmszNWIoFnkgBut1VrJaCTfq7lhF1H0Pe0zWKHcWBErW2XyRUjDm8goi+
7lAyVlwqeVHBrBklJzJ+9n8euBmmdzxBXLs9pXaXvkmn6tnYZ0g1UTemfsSTqzf2
/RQQUu0HaapdJnj4m8CeOuBxThmYbjZuHvKBa074MnajjZiAZYB/N7pkUiRJL8lq
waF4aTGD+1uLNE0u9N5LagYkvx0yvzTO67D/O4N8wP5A8ybGOkvdOxDfZJ9rfADw
FuwnPhH9LhqB7z+1Jx4ejy1+2dgSTOnrK9sQx3J4mSsnXQg4oqxoVqClavrMTnia
KOcG0SEzDKzb+pN7Fzw4V+DV424mSfBEg9TksaxgDAsezeaYhmStUDJK+1tZTgYi
HVUNrcoU6f8RqrXGE6prPDKPZvv08kNGH9dEwm3rY0Cy9uRwqmVN6lZNL1rMQ6AP
D8J2sUITo/68D3rJ7hNiZcNH4nwtV7DShbRj4jGN3xpA4spM39zY5pE7X42i54DZ
lFUNnlHCRB3euRdYTm8//HY/MyKuPJd0KrTr598LGnOfSPywX7udNI2qZgZwBBnc
4/dq7q3yETL2BzAxGZ8yArUhoRjUMNXG7w7BoT4PRT9NVhrXxobXhxHJ+tPoASRS
ObmavVCl9xO5i/8u+PLLFzrerTorS4MsHibcVyiIfsoYZNeL87QfDtPMQ9VhWVlc
nJCT29OGFxAVlQqJuK9FyeM94qQ+pCniEBrJuM9EJZ4R/e8VtX5WBo27/pI6fZKn
e//MJ8MpT+jqS8AagywY4wC4YJYaBHxFfrrhvBO50P6NiDqTgBnfU05PVe6X13o2
0Uu2uwfLM1zxl3gNxnyDefOulPd7Qina0LqdCyX66g5PmkQvIuFl368yaGCfAvYD
jXliguwhH4GP9D8hAea0eKvMz+JPnGCR98kpd0uXwhI9tZueWMQDxMjGYifWJgSi
hzerEJHWc8xOpmBy/CGWwy1FeVchKzvxpCiSltx8GbmlbFvZG3mQkAHAdh5leTGu
uNbX0lYBoq/6yunIn7E4ePIeWryv8TlX27nxrz+kyLnV+3Ahr7JLZ3g9n3SPkFYA
jTdivImRBaKsN+AtvM12Tmp/KycBHMwICm0FECQXCZkgMNQf3i31qzE+P0qnVqLK
p5gC2VJMMtOP8MkwrK8UNBQ73FCdjVY5fCBbfB0xNt4k2U1OePwqaIhvimLjdyTH
SozmG7vls7LHks103ZvEA/RQ7AitYK2bCIwUmCZKD/jUs/UcTaQiWFje1Vkdcccg
XhMy8YzU943udgY2sD44TYca4tuT/McUyPTlWxgG3oH0WmXAFVGxrBM4wtuQMmsy
s1nXVKeC2AFVhVlmDLtrEOjLre7RG4bGxrkTogEz9ZYDKpsPplTAGvy08pWVI1Wn
MKfgRTm7E+AToDvs4e/gnqm+XRSBi3Yf3AiKCl0vorOP0Tf8ZfkosmjK4P4wS3/S
M13VUu4Yb2kEbSgFTlcv/uosSdQcS6x6NClyb1V4PG7A17gvLter8HXj6upFsQvc
WbpzdPaKk1mXjjREAIgTdKnAIAlNpgLyO0l+NmkJsT/hZoNTThOLbKVeLKKwlvYw
jj5cuQPwT0LBNxXMO9UQSx1GrbVnIks4mQfDUU5I3P6yYDLQlsNH4GZEdvImRbL+
XcnQW6aTEpB5xh1hG25BRyw05XVNwIQlpCyvJb8YzrLYNpXJvEAeh6DXH2HfFwMu
i5F6P3S8DUvkns2/O1xKj4qZ0/mIPPl8ZfEb+qWjaW5lvnGAZDAaJ5cnOPppaHs6
BjF+VsxZ9j0JR9TNhOGf5xmkyuPWCbx541lvFLhLJtNN0l2h5yhVJeHgBD/d7SKH
8H/0AHN42MnddkS8qsbO1BMeUZmD2mkHO/HgD3kgYv0eZeN5AUAf+IbpsS9yTSgm
jGZawzLyBUahyaQf6pvkE8eagYHDukr3fOJHvzDZcwwQJdGc+X50VocPZGhtaq7a
kuzGvFR9plEnkAA0gX6taeB07NDDuNn7b8jGIf6MDsg9iYAizGaOrLDnxhKxP8Qr
YrubCPpXY//gq6qAFYO7Chm5ECCh/5BavoIB9OQc0fvhwsdqdKYUY6PH0go9+J1+
dHigH6yoXHnWxe3wifiPlRHo0OWrUKMSWNs0wTE23AxH6N/oOAZvW2nMoQsXdFXc
eHKOH1P0MdzH1DhoM5nVQDKQHccq+XqzCx8/deYFZ4NlzGgH5PkO8PFoM9VmBVLV
YXbIdcFst8dKQCtX3xB9N4pUYEq1EgG7WSX20ESCZjJGz5VOM3RHSKv5CpUXI9mN
GE9rzKbVY2dQwM9obGGO8F+ChYMNBEs8u/ISYcUL8BJhibE94JTBdcxNiW7472H5
QFBDMOfjlVUxj3MHQVrny8sz9y/HM006HsEIJuuLTVHHp23i2cHWIor2uQD0mD4V
KA2N1BLao6GqwjtvnNb5HSh+jY/2DAC3nAuiAu74Wz8Jagp2Sm4OY2nD732bd3Q/
6nkRkvFhTE/sI+2NODn6H5IrDAeOjc+VYFQO8d5nFb7q9HaohbpJM8/CdOzVQLDy
batzuGkRkuzkycjFVa+HAxUqbHBI0+VbLNFt8Dvb1BzJcnsJ7u+eICoZkcnTv1KV
zS/FxVdkFWqkl9VIoLs3qdi8HrOlgk/KMJ6NmMQZ2cvPbV1wJjCaFFV9U1raen52
YHvTQ9zmA3JdLndDftflW6wVCtZEsoGpvmbjbsGvhirCoK4GEddozyKOUicSofJl
XDmGj11dzKd+w9VnNOWGtS5AgSmauU6ChC/xGtlSaJyMvkzCq9D0z9dJ5+rcO2wm
am+Mz7JQcvLEsXiLvhpFeF9PSE3z6gUgTTJTDBjm8ohoXF3KIocuBHSP/hrb4D5z
SCLZVMEKm/uNVEt0fiBz2Axjd0GXKvFFqRCOmgK2THk/XWAGduPwJf5UAeVCU8tk
enaU40R0oNpw2neO560/Q1aRYgDUdJlJdnyXDs2rRIID78/AlvzQpGTut1UnARfH
plRvB1pdkK4a9GFbT+4JKZcuxjRJIj84En1uPrkVyOpGNULHKwLI73nS4RQnx41W
3ZkunQIgZsGU7qQWZEsmsxF+J8Lbi4fg1gMwzvVtbtmGjrjpTzQkIg5HBdoQr1zc
1sriRHMlOU6jj83uQ437xU9lHXXQXby2q7+V0yBbIEr0Sgjc6RgQW+1IUVzaYDA7
akzvOdU+WiaYoskJMmoitoRQ7YMMmaKiWj08rA7Pv+jwGlSEJ+N2qNR80evpEebD
ptGpURUh49VKrMFpBB7UgwYw7j/gp798BoLgBdPvjHbm7WqGmU7jw/NeMrSrt/bJ
sNbQ8kux52XNJBzPVaiFjRgmKeM4B0QM7na3KW+JZIQLIeK8lMrzFE70IrJtehfF
coC5qCQo/X9h7/MpdDpgPxsWXqTyJLiTjIJ39PY9N7AhojoSqmS5aahNERA/eXmj
an93as009Fki5wK/BtFe+gJEfXhn8k/NkVE+pHPK4kCquVJZCh1jN+m4bzXZxyya
/CUNt8WbIm526BAYbE0MZHVJ7IOmJDv8eo4ygKdp1axG6GRgOV/sAgJr82nVN8fT
mNPG5/lTC06Li6fKfu0DwWlz3M0XzmOLAA1sEtfXi3erW0878BWhTd8azmQNK1O3
iWlfy3sHF4im4vRUyuWOtwzhUcECNxKCYWL4bjQi/d9BN9IRNDnAD3Q2mQvmcp+s
uCVpPmb7nXpNfmTp7n/PzadnqWBbCPxmKwand438Jg5WiksO9CwwDLW0mCjmSDC9
w8Kv+G9TdUwNfgqe+rxh0oCoMSICQJqeWrrsLuwwKElFQ4ftra/WBaNiyThYWbfg
arabiQG/OVxikwsMonkQCDHA80Phoe/m2VYTOqJUWbWTBiUWlKUJVqYe1HJlknl8
+uG22gihWQ/zn5ihPLMSvl9zmeumXHK/w28/kKavSH42PFQ/QE4uBDrwYkoTX2FO
JfEoNZvKwZ2gJ9/29xoEumMghi5mcYAQPEC2SCOginzXVSq56dEmPP+o76bn+FEf
Tt51DBZ3jn7nYSGydOEUUPBF7bKFLJabpK7lr2cDE8lpEG8PGzYxSGVgCy5RDVbY
XiOMjhWJ0NDxyeg5b0+OdxgWjvpXAXeihj0JPMfF5LacoxvPLi//LBU+MHHSTpRi
fEYB8PPR4UASvMiYbH45fFv0nKwSqa8WK5Ylgn+ClCxNEkr7PeBD2txh4KjktKzD
o5fvsYpPHGNrW0OX6LupBIndJHcc8SgjlOjRBMrk/W8SoktQvFkszecvU0JavGsE
hRy/r0MfjNUAaD9LCkTKO1ll/LWyn3f6zjOuErxam0H5CUuIKqSsln2XJCwjH4DV
8UJr+K+qj8gLr6SFGvoJZFNkKaHXzxe/52ASAMDN5Rv2x6JbGJhyXhAqSts/crYK
BTUtsZRabKLB5GUEpOwEVQIwsQl3mUACKU+RgSAko/IDB+cFzo+WbWTVG6YT/i5B
iq0kBoAblE7g7sC1MndInQ1sTpRhUjHsLrkZbiENiwOq+jphXRPs1qGKB5xsEXPB
rF77MwQ6AVryrkgcLjKOqCsI9E3WlLZD4Cy4Vjnq2HGwxpHIPcdCyTf3pmZwtb4X
ACSsvozx6Z5LQyzfdDEJARGV/QItzoOOvyb9tlRiXE9dekaTbb3o350B3fpQs2LQ
lokhWH1A/mtKZMoHlTFvBgPL5bJr493X+glplRIK4oC1Er2GFUaUPjgyvkzLc1Hz
10uu2i/HyoHxWeaIpaG8GaXJO0a+26qN5WDlhXcWzaZv2mFJkeqf78oWnr9iK1Tt
vkn3ZGoo15tZGjh9gFO3sa93l3sh15j2kBdG07VDPlxLzFv8vDf5Cn30fQcbRAZ4
msLEAX+wIsGAgX1en3pKUJBXZYg8S8dZVGKX+Oytk89+MRmyc7EdjqOReMnaw33U
Z8GQ8wxgvJSVEhwd4bQd/Eyz3aAC1hvwLspYO2TL7YAjUIoViZrRE3215GcayNG+
g1QQqqkorcoX02HV6AJ+uSFKLjM1bi8x+JgB/MmLkwkU+QTJzOFZ1KcNjgnBsqGd
gKJbIdqVVRnW6Ps7k4a140mYnAzNBaWN5hH7IyHEul7bOap4m6CD8PUNGpTCkSfD
AJI8kv3r7Vx9z+o4b8OPUCjDWTFSOU2XwaT3tJRTFHNGJoSiS102s6zkC6pWAcpR
hPzDi6sndYlcBwTCkrUHn9bj2J8dVKQOkJziOCxcsZvtIXP4FNZ/3487V1RXZkfT
pBUXmmQ79Jqu049V0xtWrpHt6YXnojS7qYqzYOCjRzqw9U63ND9zicrXMuQZTpFC
rIC+U9s8QmKZE8fTzrSC3AjNaqnpVk/wTA3h+CTUjyIrkJe4Ns/CoND/0xa0iTbj
ftPhoSHPOIpUBafI5KmnQRFp4tgc2eNWcmN18jguwVJPmWPNfTzgabw/xiamNgGC
Book+RSslDS5h5Go6uHjY6POdfVdzXbeeHhS+azeD4U4yciw+97Hwvo+lFOzbr/L
/q/gcSs3HzOHiw+guE5FAi/61NG03DzSFbyle3Rq6AUQBLgxq+HRGKfSTdKtzn9L
2zv7kS+gwOxKdyT2FAyU8NSt31cvArxda/Y372X6MUgyYpZjC2fH39qy58BDt33y
pZDeh1i/KZ6gPCAqlinrCc7CYFbebBDKTvSH1c2ykEDByUCpbwEuv4NXCJHnrRXD
XrGXU0qepdqRfnhfB6bb4YstQDjfjBNJHVLLW5LG9Aydj/QZWM8gpz9iK0tem3/A
JS+Q3jtcB44ovTzpFNBaXpsihqtxMuZkLNfJMNUhUENXp5O9rCNS46di+6u3r7T+
C3EHBaqW3m27IyWQ5XdqKJ3vSiHzRNexFw/LubcGojk5ihU91b8bfIJLjKoNU2ps
o+0zd9jgeZw+6du7ggcY/E3+zY5xtYxRQMow1dR4ti3dlraaqLntLXAIYcPdKTOV
rfHWSi5DleKH1ntNLvNv9l9JLrmEzJSlKc2iuOn5tC758dGc7xV34WyocjxVa3Gj
W3tPCj3UyM5KhRZSGu93cohmr5l2ezyPZJVWjoQxBRCbNSejGeAx+aAsGoBADDkl
MDNWb8nxtMJ2ezcZDbDH9YfT5L/qDjLOOw+e81MBsvt8fo1Mm3bC6T6+0xPHEha2
TDieZanVNPqT4zNKUt6LyUhKyeBaK2bBf7BXkDyuvQqMXHYQkf20jP7sMVJ8K706
S/U6Ngih0RPeYzREx2mj3bH0DEH3eI9pvFpzPSnTodOyI1SFAEvxhCB1ipR7dy0o
OncAKBWMD7KVWSiHEVYLvWtnt5Qn1KmFAQkDEns+wZjpDAieDzmrD5Uz3AsVihDq
ng3Z7km2tS+/4OJDF2JC2SSj4OJTvr+cTKHJjjjw98qUCCXhjAvOOgU5cfIEorFP
JqqjamATfKBOT7hUtSLalTehu2kOhu4pGTulyFJIxnkmOiE7nOJQvsQrAw5XkVp5
a0Ih/t96uIl/vPKPRUkubj0MgZsTX718Au5YsGL+E2K2nE1pvaxi6/x6NHGtrlB6
ycvzIZTD7zeVQh27D8gEtcqjSCWqoENpdnXcj48+Skas9vAHyyRE3eZ8JAO7/dYa
uM0l7uMppXIhO8/iaPEsWPPm1BJO1e/T9S8aF9OeDOqaYRUR3anWfLK8E7Ir7Nw6
CRkA8B9W1NB5O/PeElRd168ueBB78mWQLV0sdckFT9Wa3UTiWnc7IBcoIw83YJRW
hzAHXVzeHuy7BuNO67YLSZTy+Bj2SKDjIi/wTiRUvg6cP4rICQp4Ma/3Gcuksyei
iIOJNKSADWfuT8zw0vGhfl4E0cfpmUwo950FoVfTZ8n8IDiHQEriPG2JUg3GXDqg
OUZnJOJ5v+2NL4uf3pPScB4CKi0KCvv4L1S0npSRYMH2ZBMnu32aRnkqvrw8BC56
2xkSzxBxvbjaEG350z9KzI2wNaCvVnCqeGloUV5WK0Tswfu9i33tc9O5Bb/6Z88B
t6ucw12f/W/4lyhZlalK+cwlak+Ghrp1rP+MIQrvOOxmpnOUD4rFGbgSYocoy+Mx
kswEb+Qirrrcla2riZmkAEc1ZIZuJUsYhn8rYw5i45qFQ7VkHgPr4TcAXQN4GoO+
ZBjDcV/3mMlpolyQ9BeZ8LwOL23BDaBLbrnljItlOpfxMXAilG8G0Y3czHa62TCq
U0L4zqBxjFEiroYH9ScFRqms+DgvN6V40vKPD3zAYTUnG7aPfgeU9OuObC6uXMHt
l2R0nhWUN6VQB34unshfEJrSjrTQMprGMfufulGhNvPn1hcO2KpItRGE+nefCEJi
qNHSS47c8pHVFg/2ow0RQ4Fe73IpWIhMM6H9pAqVs1vaXxdk3BHCLpYaGmbAo236
fdz5EuPuql3Zm/gamAWpRSkdhqLlvt2T5P2iWddgMIncjfAvB1U5i2awRYzZm1O1
WLLMjLcPkSmr5Zc2knhXFuZfJAIF/pPyHQRiMFW4TtEj0h1HBqItcfXMiMZVSExz
+j5/qXbxXL64LJX+Q2iFFn9mrlUfkHG0hoS7WTt+HvR6YF8HgbGtX0O6xqz7mA31
UJe20VI4lXopDLYF0CKyedyAho+FnCmyW2ruBjQgqVWCfmS8WKjHUZfq3lZOLvRA
6LNcdJHxW9lZE/eFeFyZ/NudvLyRfH0eaVUGxlCSbuMfQvQJdV36j6NHs16c9gpR
6D4BDeha/zjjo9dtn3hkLiXNHUFOJJgihcJzYbNHCDSy94wq9zndmrPk3e7TDN8X
2HousVFVYAm717yVvMbzIwjkrvGKc8gNy9fCL5C8F8BlHeqfdLNMMZ/syHfrRNJz
VDqN+q/3rSYsUwY5kVlKmrfthhNMGo+kftateZeZkHA+0buV6wrhz37vKVI40RYU
mb0oqfFb8+9vVXpfCwhVEDM+pkR3Q0q3FkeKl2bsJiPHB7b2Kl8GuBeZdUFDXfRV
M01KL56ucBztix74Ub0CQAUafvLMtiuDWAvcv5bRBWTWBX3ljGF4oB2nts+3VdMQ
O4JdsuKg76r6CmJrNy4XT59I+tkQX7fnaVsVkXsIJ6XlcGBRDzpeXn2Bq8CpQfnW
0CbziY3WZqwHmTBURB/++wDGP6Wty55Agz9UXhUDUDvLDpiTDTxbAidc1U4jsTYa
hfH00qCji4ATmVJSfgk/QbKha3dy7Vn1EJjpatXo94vIUUQ49mKLNxUpokzaYUTo
LC/M9kqnoO3+UJjfje3SLBpEt6CD5mFCX6x+s44CRkPUVTLwbTD6JqsFjnjb294c
te8Lh4gk6xgU9xmZUYT0FVoRj9I34Kv9mdEIiSmFXoD+RdHkU72KGnMMnMBYQTjh
oPM3gAa9h6wXeEFnIfcQHryALQJ0gNVJeRd6IqFpliEJcL6a6vnbqJZ62g8cFJnE
yrQ69MspEB7FDaUi9994mdjSZxw7Ms0O0FXKbJd6XK9iMp5Fkgz5an8ifo/PoRrF
IVTtW+YwpCNsYyE5B4yduTLHV9uQLv6brLsrDnv2JTCCHXNxhANkNFRDfi+ViKTZ
XCNKLYXENihxBeepq5O1iyaLamZtiPN32ozhoq+z5EdsqO/035QGEFW7rXFiOVoo
10WaJaKHhwqhcg2MA9Pvcypp5QIIOgOQJ4Rt6WRhMilDHO0d+LN/oeOmjxs7R2B2
HawnN/bwchQFnB4pDNCADErah8ONnLSkvndr99BgpkbT2K0333oryTLiwMMgvENA
CSuVRfx41RgWXDSX+eQFsOR8XHGqerOYFUV29CvW7Gm0+LVybC/fhDTVi/FxGQly
3iz6XeeMzNORz1RRyjmRdZ29jUM+FHG+AvtS13yDVtJ+/HP5NfcyNQxNiB1Ckqtk
8e4LR+B2jFAkJHcQVVff/dC2VWaqQ9WRFgKzSw1YW0SIySl5pS5ir8fCYcQSPCe+
kQGdTzELzkUiKQVa6L2KL4U+zVJyfOfqORxKFHAjO/nfhH9QSUUyaKYe4apjbdRo
4DOh86DxL1F+cmAwYAGPV62m0EAzfhItXR+b/Dbm8LQIVeAP5a9evkC5HTEJWdUl
n0C+P66KBSqZJGhnCaysEYyVPVkEq+3qlRRpauon+T7PkqWfyeSG+Y9O621Qjlar
86zKwRB3GD1smOWfCjLaC0GlQq2nGzyBTFo8Zy855GK4uF8T2mpz9ex3yyMILAgE
OIjtCO3gywubo7i5Da83mM1b1JqBPt4xYWNCkAEQqX6eq9lpk8dLCliXe409oDn6
qfdBaDiduWlwaPbpVURD+dvUZEbV3pfIxpadvmA8jJJinfbgTLgKL3/s9CFl58Yr
sSYuxNL2ow1w5DQ8MfwNPJ92S2BVxoGnkBmeM0ZUMZk2OdfOuELzjbwMjns28zaa
wU9Zz4eaXOd/zqGU/iNaXji0K0iK3I7XxiWS8XsCKYZ5jZHDP4kn0edPOSjcMgpV
UcAh399Ym8EQLZqSVCsMfazvSwZKywjao6c7VIerXCQPzGqF28+bWlxSgDiXAYgF
iPtxtuelBn0qfgypnmvEEuunAW/gUcbm8+NA119IKZ0ThPkIYO1u1zcm41njBjup
r7FrR+8aoMF68IfVnWhiT72w7aNptgCdWOiTE88Adq0DImHvKSo71sq2Pt/XR7b2
8O19OKp58UorQhGy/gOu8H9aMVZ7h072i5hftsJKzY84YizSsHIbC23kevpD4tT/
r5H13OPb1Y3hoJeeNrnYPvNRMQ9NP0U/rWazp8Z0M0zyXQlkr/UiD23ICskS1LwH
clyAA5wD5cAhgzYes2JJjIwYTFUG1PDX6R0xI/BfFvaC0QZ3y0STCqYJLd6TZoS0
t7Aa41AJPo+i9PuelWFKpdyWiJP7lb4a+GhzEvXUEUbCWZkaP3QJzMw5fKnwGJSe
V7pwdC5fRosieBGt8yKhJuxI7N0EOnw6goXSQig2Z6F1K8iOeB34HDPjJsLNryfl
0uiodG9+s0vootxnPFjShQoT5tV1zgc7g6eutbU3JJ6rO0t1O2sVOnvK7t9+56k6
pgKwyUfR/BjmJJf/QKS5x9jnsJoeYD8sol93ywcrHjC6gKrMQGY5WNIFhUle3OjI
+aVVxefQlIo1MGgUB2SWWp/vQAYXdsfTlww4IO9dhFuw2f15rbJHw17XFlhHVrm9
zKKB4xbkWmTDFz79OVSIm232jzWZd07XvF7RNl2H77vCJ7kOr2ffo7nHH3G/f3oQ
gQ+LGJMD7tEhTWb42fD5EoKDsPjyyR6QVRmNwuLHxBvnyzVLuzif2PWRWOXCTPZ3
7f6gs9Pd7Aep7EflGxqOsSEgM+yLdVcH7+dmfUKSFjDr8MQ41LCTLLD6tPHvO1+i
X/KwXadh9G3UnvFD8Pd+EEv2RNPWUxygcyoIV225wOlj8RR2sTXM2Owcj6hstCw6
a2gVUizRivPvtX1c6KdgNWQudLLDxHuGkH1e9Q9i6bxzFR+VCCkh0iATgC7X6Z/R
F2twcA8O4jAWLV9jtAXT+1OBaamovGZt7CNlJCw2CwctUJCR+cBxLA8AWK/0K7rG
Mde/V3Mr4ZezQ+NsiK/3MfEcx3HJC0PrIVwbqNlS8rOBaeaDnXsHzfEwZNadnQrr
AajoO+WFSq1dzFaCSY4WhadYKLt3QBIrSlYlVY31dcU3RfeoLAy0z3DBo1ujcf1+
UNgs3J/yj3ImQOry7ucIEEc2j0c0q+/QXp9FBYMkBAObsbzxQHAvIId7Aj1RBJVR
HqCQw100HzjOTC/V/wLy8oCMaPY4kruM9yrjd0M5biZoJ6lTM7MnEdgI4lwBpqxM
Ianlx9VR9K3y04f5vyj5Fh30U2nQLT9mxvcg/KRTVVL0xnhqes72JvnDb32AXC+p
MR6aBNkmx0vNdcmhvZCFtdsiSqIFxEuTIqnkGtn8T9ir1MHNyjtdvd6zD+VpoHE/
QnY0S/ge/9z849cRjXYaZM4G5P2hEZ855rN4R/0JmxT38mpdURZxM25ErxTidCdM
iKwq+X/ZF8mptO9eD4ds2sN/cl3Qw4tLmIgoALrqyvM0AU4f4PskTkilmGkBVjyk
Q1t++uu1Z9984deZ6U+V9jMjn3PFd0RRyZJ4mJTXqEFMu3LH6V/Tx5w8IVZAt355
cxa0/xEF4TAiT9TX3R+qIpHZHguUWQfDjoeHwRX0tIIT5E4NcnWxv2GowOzM/vuG
Mj3+vPOHZs7MYIyxANzbsBjhZhD76krLhkers+RfL5Uy0LE4OFHFqEcq6lklX76e
whPqSvdLvvdmam9U/NuNsEGtqGhlXSGJ0ZiIguvBf4HB6SUgTxpVYhmrInh3QMJ7
pn9xCU4NPdlnHtANC3afemnsX9uRM/m3Rh1TKAccIvZ+RhcLXeT4dO5nHR0i5dy8
esgltALKuz5kzOedZeybj4PzlVIQprXpEn3MqsFWq0rQFabyJHkk31c4cXG2df5X
tfoXxfM8oxoiE7fRMmOa4UBQdIrndLUO7fSzYegdESMVnrabLStHZnVqnBi0HIQ/
iusTmR0oMk9Yu4RuBYPignJylPYqU9oIlP5zCpN1RmgxdbCyvGvwVkPyhRuDIgGw
nxiwnykDucskP8KoC3TKWke0NhQEi9rCwCBRWM8NJynGnam7Qf+ImICv9xzxM/ik
22kR/pKAh5Du/nnV0VHmDwyEaBX9AeSnLBKHRPonSoB0ZUb2mt91xyeVVBAhfHVL
sUWekQ1529MScUOMjNb8iUOgH/xR6Z161d3FA06jnInP+Kp37Lgv/DSxXTq4YBS1
M5MsnisWSNFpxR/5uyJPwjpYz1K7SJ1CCoHRw/9wO1kXgaIHXg3nhcSX5VQsd0QV
5k6OFVzYUIwue/57QZrvUU094gMeDKTAqaSjKf5i+MiEsqEmFzH8hl1V0tHmUqHb
s+uPteJnIyGz1yNyp9DimQUlxrpj9hAwyKxKvJB1ZoXVCtPXzlbgABwCfjfjNVTD
9v+ppKxr9eXUa8hOUgvJxaSW2Vv9W21F8zwFUtNLNOa+kYNhOgQxvnUcIzxghuKc
WA+ZrxvbF+HO3q3CgXozi0YTd3FFVnQZ4pKmuve3zAPtW/4WI9Yt406zpJaLV5lc
MWzQQTTMK2tQPzcHOByhHSDVWDToO7ZrDttrv4Eqtke84usfPvxKC0IMMG53QWwr
0Klqjx+QVhOgggz7NaNcWplhevZaziwg4JktDGSrU3WK8U0QjWsTaWQ2f1Q0PUZN
w+/xkULXrTai73DhNkZDL317TxF/+J3RM8FHgUshakOchlCr/Or6ROaT7KgpkdTp
iYNFcAcq2ynihjyKg5MmQelnmzaRR+NCH5AsfMSXJ3M6cSon3got+c/rHAMZ/zNu
AB4g74VTb2Vc+iLndTnigBJqD/ncs3Kn+FKEyqPsHTNcwDx5pFIr+gqr58PT4KDF
GiPqlhy0/2OT2T9L3ckc67QEyKWwll8QmD5hwisxgSQwpYlysP3aOySw9fV37KiG
qwbvxTD6j06ADLxh3hQk7QWZ/wFAwbejjQdmeuxBIPFDgvaCFYKTDRxllFiqcPcY
MroxyFf/wiETUM+2uT5HfYieQ3UXJy0P7b5bj52R3k5gslMzbV4vfAvBqBO9Cfy9
Gn4iiCz9wDnNIEHqJ7s4GSUlzdfIdsqMhp9jVswlkBzqMuaotO/PtOhVGdm52Hq2
lH4BZrOj0uyxvxryeJM5yS3bgmB4TWsdGRpvF0mgZceBuNyRUbdnDviiNdMDCz5I
M/yt222Xig5xh5+YVCRuLt/n8baZ3RNEtXmrVJYln+5+Tp+ulV7okRUEHp8v4RHA
OFIGJaMCzbdGrHb+eMQ5HCJT8zxq8hZJxjAJDtvhJRAgeaBekO3ZNXRp2XUDzxxg
dcsOFCY2JLK06uMnVFvyknO+dlU4ql/CWvo9aKxk6d5Te/gGPv1bGVqftVIDdKCh
bqyMQNOxfO11o97EaJg5JNEFjXgf7JDZb+Bp80lIxCWRUYz03uW2MxGvKvQ8iBuI
8N2b+7pxUDmFb+ypl0bqCntCg8Md/qtCP0voLfiT6Qh/czUTkul3iZnlo14oUURH
twmFtRAca33HdezSMqXm3gmpewttKRLQEZm783m9y704KRIShhhDr6cZTUk7o9OP
hUKIr8I9Pz6WGxQOdwcYTaCA06gncFqzDfO8W93DzWyzDSLUQ8sCyFaRM9iseceA
qkADnqmAtOHGlBHCdAHZM/iYmDY8roO3syZl0P/tczLeCk5Kip3CZcMK5KS5YIhr
7nqML2Q4pQjVy8yMJIgZ5aDbNwArPllg3kkZW2omu85SDQe/ruHF0YtLCabXviKw
yvkOB9R/986Y56fdxhFM2xfo4HuBAK24w4yQeOY9P9Wu8OOuFnLjQxbUs+SQLSU/
UW8evDzKDtr9gYm0PYlis7zcspubsEzK/cZWlhNl7k1se6WYu3KX1FOoqG5W+SQM
yTBsbvORJvBMd1AWit+2PhjHBxtwXw8/RS7Sc3+GAc5MGAr5lNiTLsDxudCIsWk2
47VuYMumLfeEpEcEd7AkqDEwfgG6QcjKdzW/LsZdTb+c7GxsitqApwQvz096ViyF
5Hc/C4NSQB+fZxM/zLGkEJo2zbiOsOFHmm10ZrBsClxKbLXa6XYyNXWLHTt4hMrr
HHSh87/iFTLwNTKNNIZBS5VkXfxGydTGnWOXkWydt/YbiFjlMmT8BIMgxYPKROPV
qkjwbLlbuyIyRxPwW9E5jSL/0mtiBROguxmdcCeEQzMVDG+fKsYnzwY1MCFHTtYv
VTldykLbO1Pj7BeWVhDj3fkmB2tH3ilGEbvM+4HM3FjcEzrSiCCv4uUUM1EJCpNB
k6/s4v+Fxuo34B4h9RKt7LHI47pTqx7uqlV0XZP+sc9lQs7AeMX2jHWaVz/Nt98X
H6h2eT7XWXYmk0n58kvi/nTStdX4Tes9+4ax7Itr1tT7MmVsTakweJoKc0f4Le3N
S4g0B/6OXh8DwCj5NMvFH1IulEDZ8TKXjrYviAG3R/hCq1lmlMZp9OlW7nY9PDoE
U7/wP8pOJr+LKCaTy6GGtfTY+YeT+NxqYn3cfd2Ub70m/b2OxnUGN0eM2GMaNVjp
6KTSc3p8iBpVVNIl2sxWKsqR2ao/2iGRU5tv9C4aIqmLTsWsg42s0BHPU/OnnYcV
KPhfmYh0cc1dVTVEp5ySnHB33BsVjUknyTI+rTR5ChVl2ZXIIk4ncirxoy35kFV7
3TfntIK4fX5XGAps+8gqq4ZwICuWQg4ZnpGJNIzVbu2Hmn+2G/Z/I76imcy1qiA3
w/cbXf4oREeuZlWc0r70I73EXnrUqdbKBMeZM8SoQgj1gVnybL+Fk78WU8b5b0Ob
n1rdEtQkayK29VBGJsXdfFiR7kQYU+d705IOOk54qa3ZHICM96lE8fT9fMG1uswQ
yJQzOeiO6tpdjEzgXlZeogghyKKKljXF4n1W9R6cfc7/vdRHVArw0t87Hs7PAEHO
o2ZsN/SJUDV2bDVlvn1SoL9OvhIEBWsrLIbZh3Emanoh8evq5JMx3ixdvOn5fv+u
ODXzihQk6qaYJbz/hANXzVV2mOptqQTediR25+Kfp7yW3+umWcFXJzpW27mhvNAD
zesmpiYsAOZ6El50NyvAyuD3aSkP3BephjOHeq2QcXeMwGcnsDkFY10dYLwYrVWN
02qUJZ5q77bgBgAGVg7ZoWwvb0TPCrPqnkAVIrI93fCeSddVdkhPVKNHaUshU/3j
aVRZM5SCZcrzKnId+/XEg5ZKeIj+9DTAUND46xsNtHbfN/ny67CbFYZGvcupIk2O
8hOhvVoabd5byW9TybTtSu7PORgPALnxqtWXjayB1VRXg7s103ZGAoV5MH5PLVz+
UgfwqAxM4XM+XxLVIdF4pGiRiar44aUxlocqfE1owGZJgbTn4OPyo9HMgDcJ3qGg
D4R/RGgkTgnwUWHHUQfSoKHTILmaSnMhxjvTg1Z5Lrk50/uoLmz1a8aBpuXJaQDB
CWs07espgBZW+kuAVW0ackAfFSWL4RXT1grN/sSeCMw9xaqY5LqVchU2hEvZuq54
M7itq6SccsFqZJwiMjDnY0QcDptdtpZMRjP1Sw7ufeW11W3LcgAfHgTwpPELWslg
scUMzTm2WMA7BqCxsEr8Amjjbq06JLoaEw2r1rR3f1ko2nW2yU4wHAhOpkqTfF0j
b0rAR6kN3rEu/2YW6VWB5G97lrbAue3+OgnTdWXaBVxgZXjVpw6V0dt7vMHwXeYa
vxgzxDDVzYlB2e08IHTvrHkwZmHoDkkL4Labo7CZUIdptOs9qSEa5PAaoxVPzofN
vbswXMReRdMqym1r0lM98laV+/DVSQTn9AxJpHa1xG30ZZkfslIynDiVO7EQs/I6
UAf17Bs4ONkJJmHz3kAN40hjrsUQqI/5P+NWuk3p7tbe6jCqK5yBRlLSf8F6M2G8
YoKdAp/K6EzmaUwN+AI3dT+e7/uBp5VjL2GAca6W9puynaV4ozsYde2cxFX+mnk+
SqJgwfVTBruorvT4AB14/wU83VJYFE8WiWUW/UIwSLchG5t7ng8f12gKGCDA4ExI
adjEf5xkolPu2avdMvR6pIvJr2tQZjI9GFpr+8GVlLWjJ0MjPRsAOOrwyK/OuBrs
k4Jg564feuGMFD+NRFP6ZUIYO5xZ9+YxrgBdebdgfZ0nGnKz6gytrGKHT//JnABQ
3g36vcpnJjxxeIMy8ePXv3MDw/+rBYWo1QEabPe2NMAg0z4i1327EZNo/eeHEJ39
KAm2J2Jn2mJmDdBleghpddo7DcDjLcnr16xfJepHUbUPbDZi93gYZ9ZBolXVD05t
PAOvNQUWHVSC8cwkNlDiCyyCGwXlQZMD2lJgqVKm/Wbp13rGgYAdLuhkfcQxvCiD
3gbV3+LLh92JqURj08NFNxXVPXnDpefvAcKJ7dEFJ6sjX1otl2VKlrDw7anjRWOa
Oq/LkOy4LLRV6IONOTlCRcoFfAk5kPZucfEoq+KP5IxibbafLZc5ebamcsT4Kqqi
qbh9Sxr9/Ox4mQW46efc6VsRHSkDLxOqMVkb0SZFa6W/L/6QYwCUt80+wKNY6Ujt
pOs5KXTWsQWUsHP+uF9Or1/pI7Vc10rjnJu4JACYwAsRlG7dputKiOXZ4/k0aeVC
pEYoaSYkWMwkvyArCY3s6IPlBF1UpzUQL4Abd8HOFFlUIduWvvfpXKWrtCnATAfv
UsxmPR/ywhRM0foX4QEKsk/VKdhFJo2jZ5EV8JpgdtdYmky7qmMpNjt6N1UHSi8y
XctZCl7KjOq02MZQYuahaBC6Jn5mD2MohSyLNH9uYOC1OVRxbx2kDzkTDnUXS1Qf
02Mc++LMHpUI6myBwW3jviP8uYA0n4GQuM7lF1+5TV7KvRcj/D85UdMo5b3OBmVu
LA7uTHX42AkgUnaRPnPtAsnKnDR9xHvbS2aO257CWLOCdp+d0shp3RDKkxkDIcdc
HeuNfxhgOQGwmhoRNG7N+9ycEAcgIKpVorkWmSrHH0xgqu+GsaCVGTLOYzEOgdXD
EgQj6Sd1EL7PYnSwvARt1Fg7DV4VyXfO1JbkzyzLhS3KHpVH3rfLQlpTVGbwzdh5
isWt9otKSHZporLpB3qR9G2GtbBs+Qp3U+Jib9Sd9VW9XN1MJwZ6v48ubnhWKOzy
KslZ6oPmqsWoP2JdNfknFk6YaDsIQnOhadRer8KpiI0nlXlvXVCP/O11vLSivLFJ
Kq1Z4EUOy+bGNYI266s4PeSsk6rdHLoX+nLHo6tjxBVUEcRm/UQ3JkHxWglhtQZf
1Ub7sYMkGU5GSnlA/f7UB0P2bx/R+P6QWAH9oU87Wmdqypd+fJ6AMQpA3/jKkmv8
t+c4Rgsqfg00dSqPi0Yf7pIQsvrFZ/9gl5i6EmUwxGRvFfpgA/bIXB509h/9o9/F
PaAs+S2/lGHhwdzU+6dWcxYK+CW0cjGPRSdEIp/MEjN8pXU1GEEIp0fdFTk2wAWO
SERowfOMHorSHvpZNbDULqJcTDcial3cJjRmmTb47Uw/5NULuIRmcll/aKGp9aMd
Ei5EC+riDQKDEvzB1YIOsuNsEY8WuyfGn313JO/4vIL2L3y4bcAMJktH/DLWipmy
LpesnSPIT9xSoLUb+rN4BeVQoK/V5QUnmuG7fWfOFMvsk5EQp+bNgAznY0xwkYzc
byXNqgtUWtu7tzUaKpfYJSslw+2heAQhq/nGkWAGfFw0H1rXApsiYidlS/VQu5B1
gqv0Pj90Gysy9w45XDiUS2yh8Yp1Y2R+dAL9OUfvx1aH1YmjxMgnEESL69UHgFZG
XdJAW/cYe5X8Fzs/iiqHPDWN5PXkAjdkigpOePovAsoiiB2/6gpwN/50Ui8P4P1H
5BObswb4fS8c+7fZVJDRW+tnWGTpO1ExJJbSOOU98mj3HbKOxP0prcT+mpMDx6n9
Qs6XCLaP6YVbqqO7MbTtg8ZVOecHjWJg5IpZoC6/lKp+ROxLRm5UPYZDd1eik950
CcJvZ/QPCWr5LmFu+aTliVQ6NRjgIytv/JEqVQlkyddC9q0N5WN28Pgjm62AXUeg
flXk+7d/9dyJtH8z7kWI/WOQvG2/B0JUs8dVgd4r0tZzrjsE3EKNaAD9fQ5KJb8c
CS+odNtmj6Yxax5rd3Ia4z3wBcTtpzZjwNzaHAndcTXB4s3ZP6eJg7GuYcF49qOK
nUb2PqWlwVxMVwobo1W4TTjOUVh4T2nvrPIUB6dXqvKngPZiwQgdd4by9TPQFwvC
WoTs9J71GpEXmN6YnRpYuAjHYMmlHQ7uz7ei3Hs4bRQySpgbqLF8D2iolgfBuHm/
bGRfIRfQL9He1DgnU8uTKgo98ezJp/LwVEF2bIFf7ED/aUf7+x0AxkkmjzxJ1oPW
fkPvvvOE2ns5zER8BZkFEewJF5M6Db8DK7zhD8ROSMKQpBRRAWp+ohcnhAH/e9fu
2aFYhDMNzqnQTSpB7lNPlKRbRqWy4rv1Wvmkll2lu+6irge38XXV7jr3Z6aQJ4+u
HH4ulnvZeWeGKMK/CTMoAdcxd3qxeftIw8VIjhnfnQaUbt9czVEpP8VqRE3Njvg0
677c0Y3vXFyoqjWqnzBl6gpP0yzQrb3ZHGJHmWieS3jcqYwYTXM4Qzoo+I1IBlIe
vTZEQsU8VKlcmpFd3QpfMj1P4kcUbwmFKVOtxT7VeFZ1hSTque9gn/U5iEesG9fF
zBmFPQoYw0KFzF/+xyICEHCgnpdIJjcI3au2L7YVA4Q59u1N6z8MnjnHAkjbuDEA
65a5aa7fkUHnjvRE0WzoL02tzrlSeV2Q/HC19O7YjS3GUGqG0fkfcCNSo3mFqgtF
/xmkoZeyHEA4/bcvKSqwjZ2gyKpT9l5MNElYHBDhwP0EeA77iBdg0YDTlKot2L/0
h7cjbQWX4WZNrXnCHROKoW76PNTrlt5ZSpb4eUOpqmFmUEfuav0T4acbaJ8+8Dv8
Gi9UsoQsIFUVhXtSSGErTpyv1A1dLmzwlIJn0cGYwor92sqXW3l+PDn59hROYiMc
K1rx179oAVaIVqKPrd6zrOhZsj2yZWrHcJGFT2GHaXA2kee3Zqk8vYWf5AqPu7Yu
nXrYz32PlDfVLhgRyw1YsKk/BJfuUDKcZvQdkJAgMJsdxE+Squ7ykivClVOrBWwj
oavf/iOSDF2YrWLWNLr+SbBuqloXWiawoqE7NgQk2Z+xQt9ufZMkSy5VoGZ0qi8W
vrdkFIJVsF9Ow4WDiHUK56NWbCm4HSQdZUMWaBg0/1NK1NnbwXKeAdZYYM3JUrmb
bX5N7pfe0U6oV1KHGFy3l/RWRKY/m9ykf+CLdL/TSnkzOaKfBFDPkry1OvmsRjsY
olCRaoIppeHC5kbxUhevOnS6RY4h9VYCHYM5EeI7L681xSa44bhmsMZQezw3+ht0
WoTOwO4qj/xygs6wnbZfCL3AcP1KX6nG5ycr72pelHqwF29htVTvbJ8wQeVyDOUz
6Tq7zfx6eXm4DeSM4b42SIsvRc+3PbEszdEFEIq0efvVZBzbBIRTMM8AsbNV6sdz
voN5dIqkEiwYOEGpztSd4/8OkJ14K2ynUJM7PB0LXfNraeVu+Sw1HXl0yTAecbWV
JHw9Qmql59XzFkWhMnFJZJE6Z4ckq1KJ56HkBcFCBZJt8dyyjwo5qtbn9pBMXsdK
9HGKsZ2aOQTbWNuyfo2NB0RYTFWn6V9AxCgt4UaDDpYiqQb1lUVRSahhjEX4S/Cw
fK32XTBLEUmyOW0a1ct7KbngouAS8pPN+hcnIHFAfa+lnw7ng/qwBb2oqIKuKexJ
7oT9cst2q9PXGIsRXJOKS6BZiH/8At862xWo6vReSumZ8Ho44hMuS6VfRDjy+cxI
QUZjvgAhWNI9w2mWRhbl6ANLt+J3ChzR0koIq0uv8U1aLQjb/TgaDQ1yt4CBas5S
nPg+S6qlIldRyqI7e8//a9dLlcmrJfyILw7DGQt8gdN4aiatewgt2KmT74ZwKnKE
c7cmPLUFeWCQIuWuV59MQJ+KLEYbowRhHbOwGmhOtzlitjF85fIrPX2yoq64xJHk
CwJxIeKe21IftW+dRElJcnNIH9VJpmavQ5yNrFaZfHE3sNp+vDIjsT+uAjt8NoqL
Jv+FoBtGEkyU5KmzOVHPEavr9GqwvSvqQNxly4S/mAaeUd5AKDibcHPSZX1XZ1pl
dY7K8tQ6K46mBmxeOic8clqAy+VaxgDxy1wyFz3pg/3OYT68ElUAgB1N8JhKRgU2
/1TkoZKt9BGozR8e4N1KvoIX53NQu+ICXxgrAyLRZoi36FlfOaF/jRrHT+podoSp
+rfdCwPwAfRqswAM6UlXrHUFU+TKETll8HA+XqIPa5h5BX6ymY142H3+LGV7cE1H
y8YuqlmnorHymQ7t7qaE60bBL/r02a+MxTbOyG6RMkLWjtcmpYfDhsdKmeVqBQ5m
XG6UpBua5H8bpjdDD1ueiPjwBNxkriYn/zwKyIZv3fRY0EGl11SdWQBsF8JoQoZn
DH2INVEF3Yt2F+8YTjoRjQQ8m+thJ6j01aUAWUR5crvtZ9kglWKzYpY+VpgEERJk
CTKUjp7yzoP5z20dpYUlpOm81A6XOBfSvExAROBl3iISInT+0aqnMCP4NKH0cA6L
peO1QYl3fJffJg/6lzsPSTbhVQv4jVgfMuevtVcmutsY6hQjA3vVd95V/pGQxoYa
cQf0pIrDpCch4Cec1v64VUiS7IoaoGabGfOswt5Ot2jiimnex/cDoNjWtDnyiH+K
gB3is4O7+x4FIkC5CKncBOl5NknxSlL8AVidEKhCKevXZhPLNZv8+8/NvWPNuJ4d
V6hnGGVIM0xV74K4TR31ha6vgOFQsJwRUfTgLihhJ6SIHCNGnWMuDsJxEK2s7g0o
22wonHbRC6Z5tX3eErzDqNzZcjF0rPmt13gRD5wNlQVa+nb+qDChTcIAjfkZD8+3
WrKrRuNVh9VhKGA5noljYhxxF2T5CTS0vREre8T+3NsVccUXfoK2Muk8G/aWBE2n
mK+2nR+1bjUORQzw7xg6hNOuQeSManKldrizosHNwZqh5NIukznB1mtLUogjQZJH
4bITLRmajmV0YhpnxWiQnXTzQo3NQj8afW4bAlKy0TB9wE2xeDBV748H68fzfViS
VioS1YoaQEGN90cSMxcmrjq3Mbmb/vkA6ofxCVVtpbfOP7MJoXGvGrpBApjkemYc
Z08g6qSJ7632fHs/oJ9R3FlPmh/kOOrHTrhkpgva1FOo8Y6jQQA4ftW2rtFgt8vc
IFpToZN/NVoKDFitGNIx+ctxMkyE2hgks7xsvjyLKElBm1twz6EsfuuYMIlMvtwf
VP+y5c+jn18BG+0EzVo1FdicsGTtjjXyXb0eTr1oFZZbrexJP01QzUKzC1HKLWB2
SICP4ENtyAi8dJSheUvm4Y904RSSIE1Odee3DWZ69gah/Ku90bW02jtUJJlAj/VP
P09TkygZZrD0jXOqA0UnKdP44/2am23SOeZshkGuTZ8xz6CjszPoGyDHJTumtPsC
kY7/23uqnS9apyFbMMpJhTXpw5Z93UBQXcQtBHsc/H0tU+ln043hN6VjMJX433wm
lnALmeyvqkBGegJ291gGDGOi86+m2SRcfuQZhgxX5E7h9In8QP4NjqC4mC/KGvWA
fcC7M7rMWQ/R9eubB2blpkwQagOhu+IJ/BQKJl5q/mK6jaoQuWwxO7gARTxrG9e9
5/2XrUmT50uBTisLlX/V9GrWQDBSCwAL1pkAKtpHBEgfUfbqCTvyLNYZEabMob1B
w5KdCzhHLla8lXgYLDir9BahS0T1cPJ9OTD3YVU8dcCBAG+zVZXSJF12y/934kV2
DbvrLSpkzm2QjWqivadjXn+lR7dvOGRtWqQYc4gaRD3hUOI2gLA5gJwiVJTSRC7V
BBA01fcuzimvk4mtkl+Pxq9OrDLlQ6+1nbd5aU5bKqDo1HtJXvZVJw5IxH95FZc9
BKRpyQpYitr4Ochr3zT0wRI667CRe3IQihA8N+8Iw5VhlIkOKsH3qfH8QVWsxkXm
Hd0v5kmyov7P0eiVacf/E/RX3qW0wowxfCbgS5Wx+cMJOn5hIvU0hoFleiWz8g1J
h/eU1+iXE9ajZoW6NDBVWE+fEDtxjBDp8/XLm1fQ1YHZSnB8LzTfu35Zq+AxesuY
zM5ZcZuS9+W3oJqzDhCM+uckXxHXAxMumivHZ7lhVDqwyLUkE8ONz0+2TxATlqeD
DolxdEEh1Fo00oIG6c686PnvtOJf5ipqsX+rAZljTpKp4NPSS4WLF8GVdMc1+zxh
vtqMp+b0G0zb5AT70TCKEPpjXvh45U21NHLoRJxF1uo8S7SSlIIvY6vudd9J3P1S
YdImLZAIkIwMtlkRKpo5DaQrwSNgNSkavoga3443H4PD15VLX6api984GvNcbIz0
qPPp1FHoh2XXCtc+5g3ajJojuRJUL8LAw+ukgiZG7ays65CNCdliud3n1860AcQg
fnTGyVxbdgKwp2vafcZWNyPxO+yXCBiqP2bzFZIeHOBn7JGoEBT/+u6PDHt8jaDq
FPaf4sw+rpts8U0QiqsG1dm5rqmBMf3MFZqy2t1iZ0090NgvNtk7I8rLIk7lmMvz
FZo6lxarWJJDVS//dP6L9C4xFgp5GgMHrLCBO+z/qBVOUBXk/wg5MswL9s2t9eBy
icjXsjvi3B5ZMWaunI2rhvMDCiy7VwYakr97eFpwt/Tqg7xlZpMuuOfGEErPzxtF
4zrvfCTtSGqGdmCHpz9vTbwfy0A0fF1USs/cV/5CMu0lZx0CsYInZxaVxu1ut7Da
m1174g45MbOXxS4CRn8LbbYBVGo8jGgB3VIWWFjuUpSyHE6WdMHwYx5fpOfJWEBw
jPAAzb4HVRMpnSiY1r69ihYiWSSwC60WPfw8g/lZfI4RxLGaZf/nv+jXsZzr2dSt
Mf2+lC1MuJMvuGBmGeiyLRkS/R6wrofJlFgU1EObzyZ+4nwhD0Iu2ItDXWDxJAN1
7Og/tXa+A4eBJJX/BJvpUpqs1DwHPS90FccmUpPZFwx4qlza6tqzjOk8nF3aIU4i
kwBNkzCgcATv8GReORb7sJfJ8DdDCI+iy3glNxrxDolNK9jH1do23oINfJNJxe0V
vyeK0W4FOdxo/YftfxsB7Rw3JnoOT+b2LXDW/L1ZBosYX3+VEopJCrI9GETRY0G+
+7+JeGRGcekMw4sNQZ/H9MufjVUO6E4rEPmdi4Y9nOeIQaxnuTURH9f0zFQASR6p
jxvkQXSmZavQ40EZs0HntF4c1hcmieOlQSFGMp/D+5g3t64+id2CXtEJ0mZnCXeo
NqLgfi37Eq/b5ymTiHaWIrUvtzLe3az3eYmtLeT+2x7+tMGuOY9wi7nPtVrD7E7s
iN5n5Nz5NXiAtGtzXR09NPWXsaEGnLeN9jhOtB4SidAwg7G905rFDU1OX8dX63VJ
GBHEfzZgnoiIW9DY+9QfLCqOqbGrWIl0+3WjCmFk/lWrh0K9SdJ9OTBNJNneQc/+
S58D8qmjh/jdR3hIQ9q6vjHDeLeTZ4jFj4P/F3dSuyP2n4PusEJMpFBF2h3SGAAS
F7x+es+cz6jzISTvVBw18n5KTRCOHdXBI2oCv031VdSMRUWmEPWRuCgbMiG87Qbk
QKs1tlzefY02FRtUvPFVx8dDl2lejBafx20pjU6MsBj0VSaZYIOFDZlf1RTI+FX8
mnMZee6nSbDAoRYWU/twpXRRf0zJk7gbouDivNuSa3/kQ+4d0ZZsAb8907ABa1EZ
gnGAm1OH+V0n/BEUctvNr/FWuZKHWBz16WGEurle9NkOgH63Va3osur/AUiIYQDP
aLmHUgWE8Xtwk3a+ME4nJ2FCIEgGtduw9hNOx1lfIxg+exTVhvb8MdL/vO31kHL1
FyRUlP6Zr//JV5JX1uD/JZTKRS3I38UEuTUwycAZz/y3sT3psMKgbTnZ0jt3Q7hd
XvH8pjnKbIjMExbL0FQFo0LGfKFDA7rRkL7gIztK7X6YbZqsHKNbFHe9Jr+CpFYc
LpEaLjW4gl2yTNUgUYdLJ6TBylwI2bRBWgNNJUp1W3hf2JnEvr5yzR7WHnFx9QcU
5VkF/veYsEgo/J+pC96KrnWEkpOP/msR2FDffdjRaSe5+3rJFiISltbEiMpXkfe5
hxwk6bTjymJ7qcaNjJ/42Q8EeeUGrxFspfYh3x7XQ68tEyWbH3heE4XKnnVPdj9q
y7QgMZITC5kj2qbZHyA2sWwSIr5w7hg99NA/1R1fqoV7FO1GhHNW2HYUfs0q3p9B
ZX+J5olskmQbe6peijCAPipzfvgV3L4KtXmofeIR8WB/QGM3+GppACkiJHKMzs8N
eoNN+05FTWhp9Z4MpslxfGHVAY4D5veORMG8El6Msr5k/npG0iF7MRoqvnyfNs+N
p5bRWQ1o3nU0abvRk6/hNEIzu/9QLgpt3iMq7GjAQzSBMg+M102XSTZn0J9HB8nC
Up9gI6Eljiy5VIJhpm1QBA3zLR2OVQ8KgZSztnVlCBDebJk2oxFlC7EULblrDuLl
5cse9DIl6ii3r7i7ZVLE+oZ67inpqEoBt6gRyzW2WuVETwSyBHrJAMocwX8Jy0ys
CtQDVDyES1iImrQxtAtxzc6a6LkqWk1bTdxiJMXTcBJVeKgAiYmO87rOc+les/LB
j9CnWrB2dwxHfZ0KA6KvAKdj9McJkbDEdMiMncAUCQrEDrbn3GRgQ2phEO7GQGPI
NnSC2HXUMWdEb1gPc3z2OTXDzCroAfa2JpScplMCI0SzJToCKOF91A+t/8YKU8uh
qTsjEZa9GLsiQpyNQR7SEcz4KxG2ckrz7M6Soo6YkE1PD4mdUYQQKQUx1TYv7Ry7
yr1wUvs0UUmlBlNOZDtl1PTeUO8TvQp1+XMFaaT4ICZRjilbPLm+ARvMmWO65MJi
HddvXBtVuK3J/Pp6N73JcqPzZ6WSHaani8YsSTsXTqDfFqMl5yNB4j8bbSykqZOL
iSUkNxQmZmoJA0ecvF67qHIqqMFxeKumjoJRjlepbZJtHCvMtXY1aeXrXTyCxxFY
jWYVnk9exkk09N8IAtvQrUAYN5YHL2EAmzrEpqGaJN5IIOsoOqZMej4lHT4s3I9X
oT+ZfvMiZ8ua66FO0r4yxcihWUQuMRfDKYY5QAr1mrf9I09wgr+i6j8qevm+oEjK
b74UcwZzzAEdeoRuT+D6lFx+gm9uWIUvLMToGIDguSsRAlIxpl/FydZeIxxbOxUf
gv46tbNiEDszeA2jXFKoIcTpPJEuTT9YsZPtSDmIWvKDgcXVs8rz04g1YT+Epw1A
AYWiChQktoha6G4/ndA9sAyiM4iMF3cqNNB96woo6/a/0oCZ6OcGYeFTz1plnFzN
waDVkgL0mBRWTFU2rkzYFtFsEwfp84HBu5eVeghZ30HQy7danIbLKV3O7tgneZm8
iv7FEtTuHsm/qvf+VFzi6JuG2/lqbjmW3adzhlAKXGWNlAtZLVM5Q8ct4yoYyd1L
2H7eUWYwB4PH2LrP3HAy6uzHZZYfeMat4pVA4Lu3j0NCMd2SiVr5LhiftgsguzTU
sgzLY1GZxaJvqJnB7bpy1QKwEqkN03vQdgHEeV4KKqApRlQwdEY7z4+TFMLFxyLd
ZdC2QAoowqnL2moUGmO4ad+wDe2JQEDpTPlz3ajK7YMjr06bCZgS7ceD2dr/oxMz
s85JM0v8I0pKdqNt+3uUfnw4CGeqEDG2h06vlEM3H+pN3FTspumHyoz4E4SUubtf
nNKsJplIK+4/+7j16oQpib7zROdHTArrI8vIT7J5h15QOapcTIDXsXQnrCyolvUx
uTpxAccs7ZIDdybI22Z6UPCAjKkZA42bSf1Nkvzp/P6ESY+cOOG1EoDEyCd+8ljT
DaxcxdeqbzIyDVMixaInWj3tXAYagC4PkFYPV1NMJnXznf64QN93GYgG3oDYLmQp
oRXILdEqzONr7ODORATFdJ3LTHN/ofjoTjmen0hIn2Gib28YRMIVbQw6FedfUvEK
uIn/lAlQsNKB/coFLMI4wHO7bHWZEhG9XOSJxCs8y3JkvWQ37vRpjifKLtFesX+t
BWTTcsyXAGrOqRLSV7WIKvQYz/44dCHOVq71uoHGmNPqFRuNEyJsG3Joh6YtPwJy
40igWV+EundQxekEWSPk0p2whdIK3t9bbzJVpXfsUNQvWdNzqtIzbO0KH9O9QFkt
uRX4FuC6TsaQ5Jgo53R/KABpbDLYsqblz4+KKINsxrgafpufNm4obQf0vSKUGUZR
rYFabFb/FptKxeH/MPeq2/HbJ4uSkx616HmRxRG3ZhB36uIMtwM0KTR6hxCb7zpR
vhjmYfo47vJuZ5PfgLXa4ZSXqRwUkTGUv3W5u06ua1HbVuxFWvnXn8Avjoa/E8vF
icP/dbrp/kXhFaxG5NUBJWOrAXH+yjEtxvGGg7t7xlKUJKvX7/bP4NYE+b7ewFTn
zdtfvfWMVK9YA31GSxy98iiJxR1G5dz+X3OOObAfiCXV76U7Jvdueowj6TtscAsu
7q66wBYb2SsQhVTTU7e+Wko+J3TMzvqrEef2+5VOjUiIrYLfGAeyH4UtIYvH6SH+
e4PFudzfte4HjsOjSY/Gx6sRiaaP0MxyBCGMi7OqTZuD6aGnGiuRAVGC8E5imn8V
Zo3LQgc7asdRnXY/ocVEy80K603IqKil6MHdb0kohIYwNp6jFbx8OpDcSxSFc/iX
6pBHA7pj5IpDxODC4UNxnHMGN9O8ZV8bUD05hJBoUXbfHJm1FmA8uWDfgRE12KuO
Y6Sm8uU8g/VVE2sKq59VrVeC2G5J61gx2LS+22w0EHxxvISaS+aO07jofP0XxI30
AvNmfrLGPcGNL6RbJUWE5E2zU++AUK3hlBpkL3YK21Smgut2KV0PNkf9MnErYJfD
SZftOHJEPkS9bKiboWbJs/GL+x5zUdvN8CTQ0KLMCGJcI/hU6TYM62yHvNoqtfpC
9AdAvA76Hb/h4p25su/LeEdaEkO5fWkqUSjV3TobzHKuv3lxwAsd7ZURb0V/5e2a
paQsiEVh5LFD2F5Py4TQePFPiHpMuPn7Sn17M/oMLgQv7X7Lx/851s9Ap9+gSsyF
ihDbxrCQAIpThGToNzTdC0qzH8okQNHFNd4S+X+ZUCTIouBMMS/b6QZe6d2tlQHg
BPgnOuzfUNoSBbaZz0K8U1GUYX0xIG0AA2RIudxAIuCEMiYzxFRlrKtAYpPAz9yP
L+4zwYIauBItGvdfOMUhK9ypTHjmil+Fyqoi2EYfDBnTUF8DGZku+CxAJHF87Rz5
tGTQqPd3EqMHWUwW0TKYrUvbfU3IEdJnbWoVuoAUfdiDT/eRmVtxTooJdg6QhiUM
Dt36Hx7bfCn36SNo1XkypfHDST+G1dfrgn2aSemnWiDO7Lqss/Jat2wMAZJF09cU
D5evvGz2XZPxLU6fwShlyVL6PGMQAadHcWjmd1NafntZxIAGRu80aWohWGi8D6qN
C+1sy/q+Bx7GQdXBvugqr3Je+K97JWoINcB7lSBqqGmsVYsXhQoM2OaDrfpGBSmH
fg4omebvF+WgG/ETeRyRU4jc1vyBff556sPjfD8qcBhoa59LwUEhlnz57Td9loHn
fQnKeY/qpGija8y9j3E9FxaLVo8rLhTqYhOCnSukj3RGs/pN7Kndzv+l3diqxlni
Q864vg4sa/YoBjt3hZTgqKKnqM90SgXsZUrR7X4KYjlmjBXW66/WNbIjOgiAddz3
jaBcscIV0hO0IPIS/hTbRGLjjpJey9f/CX2CsYbYs6T3I0AXi7Ud9uQyU2M5dRXy
XG2DQSJjFUGkZHT/2A0TPrSbbg8Si37W/zVJ4BMwX0hdRapeZWCeR8IGHnapLw7z
lJSnmr2wZAG/xE/CuL+KuDKmQA+oW4ZvqANlhcI6P+38fXwfQUphZseubxzEAPVu
w2Jhcqp/7E/aFi/U/ZLW2iwzoovu2u9gI/Xx5ijvAMjmp5ospcY4Lk6JFfKXfB8n
HJtfma+4HzPsFqMxrtGer0rwYA2v1Ly4su3Q1QlsVJczZpah8UgPQgvvUxAcWaTh
kd1w/PSy1LXc9zr7sUQ7Fu4irbUl9pb51HuIEW786La7CMwUDV+03Q5xpOK0P/x2
TTj61pyy+M4CQ2eRNHxXu7nD0ac/JZLTQzwJY+u9d9r0t6X+1lhNnZfGIixNMpbx
IIbnBo4FcUk44VFgIfBjk+cmf4F1JiEYVkSDdrKD1f97ozBKpvAMNo38c9U3aVlp
Wfd3btYDhjgllw+bz2vJafxOUc8Fm01w8FT8ddDQ/dPkKflQ2iduvviFF/kY02s2
wqmGitan8A+TVWssr26Ha/0hn1r1CQq4Zb94WtyR59n6+D2qi7GpGueo3MywjIdq
vvrXW7kXZQ0/WCXNf1kWWC9SvAjGzcQUI1dWkm4kIRQZvO2aIgIaYpPTpxUdMEtF
EoySeT8QO2LKaH3xNgWdM0QI5xV7t8JI9B/Qfoh7h/q6s1xOpoq2fcyM+kg61/es
Xw21gS9sLGB2ns8+9UuFjv5Zr6mknlAekSAFt2mN5ALbGzb6tT+VGinT2GHgPF3j
t+8A+HQwzNMNexwc7IoYXu3gA8QHfhdJBgiKL5f3/JX/aGhUd8HbVpwFFg0Xybfo
KPdLaiyqvBOE6FLOj1RmcqUwefxkn8f+jrZKVonQA3CALwZSQgGfKfoXluZY5aV7
icTjQkk03jlsSCmP2ZPbdxeAYXEAvicdOuQ5dnQHRom8skit7ADrDmx7Cqtdj1wT
+030C0mkZWmcGsvXwb1B3qhlcVAiHMw4gEX1LYpPptC6jOfbty2JPyJqLgY5rb7n
1o4ENsqKDxjOAf2UlwNau1UDPpkeA/4t3RKMXKR3evzmnFXx8KphXnY6CS9nlRHX
ol2F28uwt07+qLjAK79U1Hze0rRqz1sW2N0nLNAtHmG74W90ZrtIFCMAmi2EjfJx
W5s9+fQODm2N1PA8+L1G2aX0VbmFJtBwY4S2yPQSSUBcLoSxIaGKmUBhciJ0stOU
QQ0l0N94pOurl8pZOJZmnPVX7larELOCmzJ62/2B3y6HMakjiHDvDOQf0OLKhK9I
AAhQPTtlkJtPgRBHgnZm+KHMjPD66r86I4EveXLCPpT6w0PBGP4xz0DrFFIM9KKm
2vw9FL3IwmpCqrWHZSsiagj4RZ8unoHOyh+4nZ5JgyuDjWpLlsKN6cotICsffnuk
voM+lUq/mzFtCNM4CenGms21rBHlukecO7GoYUIMC4BONcPeEM8nrmp7Vq5pX1vK
EJq5PFtbCJ+qevVVjJIG0VWq4qaKbtkoSK10CDgE9Dr8BJNDgTjfN/eqy78JVtE4
hAAcmI04MdnFXAshBJdHqF1vcKEif6RqHDFTGO/B42IIa1KJDvlRKpOUShYf3CbH
Fffh39ZiSyxeKTCvRvhKxSWHELifrWm87kwumeT/pcvqgJVtVnkrBZEaZbVbqnxz
BRH3Io0X2D+o3XsLzTZ/y7m5q/6muRV06+srJIteFmnaozotiedFF7kNTzShXKYO
HUZ8/KpuRB4EuW4B5n/cy1NzgfkB2c24MIPoDMVx3wIWfoqkvN7Z7osHeE4fLo4N
zYMUPDsImWrkmVxZVLKXr1MyLVEzvBLTuby7vAyg78pvrSZ/gUpu9p5nd4QdNJpt
klh1u7BNV52XGYUmdty1RwvN8wdvqp8eDO9aGdsjslD1aNFWWdHcbhtrixW7WmKn
z5LkslBA8FrDllE/ETMrD5/bSgb3QjHoarHNOD7YS6btr2xGu2FidZVtokcUpboP
ZDSG8lE3Pov6bIlXMDYhKodHKd9WHZ9LebcU120xPpAOIRrsUYybXxxhzAKH57xR
cSvIjPCeyK9wmd7SODmiXpv3hGOAgj+51brTXzLwNmZUhYJb+ETSzFPjTdk7pglt
c1ozcTQX8ZrzLhrRUX8HIHolMnPpw/yVTByzRnNj3crCDD3ARV53iR8z7RrL3hM1
P2ANymTrqD0gxAHtAAZQDujVv8ihvfLlFqSJi1/hBQuetnTMO2Tydb5TQFm2e0L0
kGud1XOtVeAVUCATcM0l+mrIYLDtXdzcrqVNcXsrrZ8gq5Z7q7pTpnirwI++ds8F
iYwhtScIVPbD78VPizLdKYgZS2/7j53+gsBOnLpJg8TQ4qLLlg7XCLrSv51w0kwi
CoMB36KA20IupzxVd1J2i+mD8jgNsJtAeYcTu+OIdCyk98M9MgGecmctlETHDcu5
HFLNBy7VDiWKyHEJnOoSjoi6zhv0Mqog7wiK2nEXK13J3FaGhBdwIEreVrhf8pNT
xYsIIOHn4h+bMkbJ/1rYVmntCK4JitekCuFK8Rgkhf5c6Nj1HZTo+9HR+f8aGl+5
C744CxdEXvw4+vMitt215P4Mvmp0A85OH7qGVRYKrZCzWpbhUBlg4UO3+Ol8R3mX
ufCAfq1cJBV4f641RfzYrQhypolJ9oIUwWyTkUKqTue0/BKfhgIPaNS3nhr2o/n3
ZWA+Zvf7ySh6vHM7xiItcHYuOZQXYx2vUaxml+Us11RStAzmZDynI9TjhmbKMvIP
JR9WyL2NAot3y/5Lw2mMq3PDe4aoZq7lpFqbfXZCQL2ZT9b2MJxvWF45Zpauz1I1
+X8P+WH2cTpW2OvxRjcDUKranayw8tA5nhbcfTixlD3JYhKkxtcf+ZftB6VHncw3
9Ar4L1QisoI0CJTDyU33+rmoGJ/4MWUyUy3W4K0Wq9pgwFs0w6kuSFtDwnWoLThx
dtZWvzcEg/tjBDnAwkM7ZSTZB/zI3Zo6crccnjvbO5BhxrP4GgzYPpsIlmB27Gva
6vi1KtE4vVjxhFDZ85bP5PVzwBO+VyPPvmoORbRmiSEeshBl+rWistOdu9Jd6sat
muyuJu/nj+ByszxDXQ5Gaw26RnzRFMLt5nCtfcxMiCa5WTDrio6Cwt2QgReRhzQ6
E+xe/3TpiKKU5Ro1ewjePodN/UzNbqmZdyMg0A3FgTbgrQimZ+DnR+eneDtBJuej
eRVFzgzHqERuyF7nQml7idQhIfNNzyrd6Yp+sSC356EI/Np/UaTHCgy+6S8Y4buR
lbPIqWRokG6Kf1al2jh9UXtOaQ+Cwos9zvMdfRwU9o3xQfZ5ng8zbk62wbl8RoKC
U/g3jFcEbTFs09G6LZMzm9jf23xkUHj6OBJa7mlcKwVDDwEnSsjPXlrcWE0p1fGg
qnEq0RkwqcZYuXrEjmfv4z0LnqS0aLO6bEOvTgxKfWx8EGVDIbrlsHXv7vmcE/hV
3Dp02k/t0Hvlb+oVsDcNrgekmUIohsA800sdd00GGJpk4liOZ5OjTLngyHiMtWgb
lXA5perfn98f6rEl9qQU8kzuWTZBx2fz8sTC/DaV9BrmgsuzjUpP3p00bVb0ycXv
mJcrnSw4jz7S4OQ6r2njO3zzGozLedzPMBjCQ9frxKk2hGlCo+eJ5ZaqnZVCVHok
D1orofSCUIQ4AucuIsb1jpuAocL5ln+V1TWpZYyyDpUgqQYrb/Qc0et/SD9ypG+K
Zb3knhe5aKKiaNqbdMbYH84Xq2rWfaqmCM5m4k9WPUASDqLZy/tQMSDOU86SpvbL
tZ83IfIFRx+abcWco90bpg3O+7EGLAralk5bc+fL9cugS6XXKekXpCS86qkJuyjI
JVzf7qnjxCXEtgVUP1YfkG2mVF21+a/JmiKsEb5rjRA+gjAo3DwAMy2X0YvQy4Fg
j8X1Cu8oqmVWRFQORoi1CFiQS2g2dJBJUzDvrG1fC2krOIo98oi+Djfjs2/n+nE/
JzI+i3eHd11BRlLrdYdsTX48tkE6E8q6enitQ1nmiyxZughroPXpOTGTJIQH8YUP
3GR8bId1FVD3JVgGoXA9Kqddaz0w1mVPgNpwt/VvQ/+jAm3BM1bNXh02P0mGEEJM
XbjBo2s/dwD4RgFASwxy0jd6vNIpw3wDRX6rQYuhLVsDtVST4qnQ50tBb98s3tZf
NpxVtjg2t27YoxbcofGWpUb/0LqdFd8Gznzqeas/NSMicN5Ax+b2zmNuCDDgmQXv
bUb2jt7ooAsPRoSPlT9JExo2oObQwzqrG8keRPVe318Y+CsDQQzCwWgsLD3cE30K
tvihSABSvdCE51nOTHumhOFbaeTGk7p1dTrHFL2VCyIOi216b6QpoaJkApDhO9qB
hhFKsTXMdJ04QLTAGp1VcReTj5c4benTshkO23SAL6bL89AtGkACNLdBTDI5mdgh
hiIu3+AdZy1/wmiRTradGIfkq6owGt9uhSskcdiKAmIAcKu8+d71VbNqMQtBD3pa
EF0buUtbWW+F18B5Jwq4hDTvI6/KAlVbADsPxqbV+STThURv/R2IiuOrNZruOsTJ
mI5Huws2B9glIHTPrbY6vWnpsaYxPXy+tJV92uyI0urys0TeTCs6d2nH9voIfVsI
ouRS0UemCGQGN3O+tTT39EOl0UyDbl/gsNrfV27ZQ4cQ+47SwRwHdHTuxSk/6xJh
XXqUdotrQfciG0Dp162p29HRV82ezV+NnqwjfQQvk+e9eRClTJH1xVLg7Lhkup1a
mM3MyRc8vtjb0itYVtwWotdn5dj8gO9X3LFcxXtmJQfsYupxrt8znSf3dtReXHmh
GwnVR8uHZEbHQvt/ftdsMBFFTxswpdeUh+DFwKwVWI5tipbxg5aZSsJD3WtXLbqa
B3UkDo7WTXNHVUdZROm8l7SXiqIXFt2huqEg9vo+zRZQkr65uQEBfcwtY7OI7W1L
fd2MEqoHKJMaY4gKPZQb9qOXSvsEy3RVtNbSdY8dezS8+djV89Sd7NJG5z6taYos
mdQrU69M6YZwrzrGKJGVTWAdByvc4c4T1WEL2uveAG6WlxJ08Qj5w1Gh9SqCY0MH
V+BcyzStuQO+kdqBdiBRvMK7BvyejUNgvvTWPWnR66wBQh5SlyIpC9alXqW48W8c
FbdOXxe4JdxbQJvSGK005f30klWUzIOR8PIRGu8Su245HA8kkzdsEuBS3rYPD1KK
7nadE/aqI9ap8ZmUFijsIKNvgycCjgXe50BZseqtsBDJDXi2LLnbLq9vfnSif8dp
yPPaeYXiLXoygTHXO87g7VWhdYrJ4291lqqRwNm+8/m1C2mbhlg+K0l+X4vLESM3
e2AMyCsftav04KCipQQPADZKf37xN59GUXHqArWt4OSWvA0LqtbJwRArVdEL2VEm
TpBX1V3C0G4Y5MOJuM/xBLe3DiAlScHWR3hav5yaR9M+IP5Qo4U7t1RDafn8b4CL
2tEbO0g6UB82u+Qsre9ZD/4X3Oq7A9AsLNs63YR1MbpGDDlKPavC4t21U8RtMv9g
/M3WVmK6RdVtEInnv82S7Gcc8jISdoQamKpKN5UZWSSctBT4g67bJgigcP5Clmmu
YYQRG/V2inVoVWMGqi0l6F/Fv6wf9hLle47hWwL5+jpVBd7HTbvOGgsNTbLyjPYm
0naoS/X0OsmGd3qE7EnDQyVMh8KHREXMLKkCORC2KC/DEZ5GiLniKdv57lOTuEmE
Nk4H4G4AM/MOg8uXukWAbpHerTFV67vDCEdgSLfjajM6TjDivnXbSX/g43oeT8DD
ExVUjHtWW81h3G/M7Sm5sbbJ85wXWGvl7igRR0SlhBmiAb92h3HVmcQOoa7nNkv4
EMVTXukFTKpNXOy4H3WIe27rlcUkbiAhBbw6KTz9jZKO7XYw3oG6kSwmlpUHC49a
O9Du8MLXVAFSkyYrcxp6+PL7i+NnnbtnJLmCGHPG4UxMF1MaguNgdgl3Wc1Dvz51
522ZLue+aD4yGE+Rl2bBCzjkIg1H68KuQa3BWeWTAo8pQf6/o9yxjqBXQPhRgBTT
VC6YB5nWJzIqWkc26alU0mq/ncB26M+8NZKugodWDhFRUYbFxB8PGYcjtwl6REnx
pYhtgN9I1kySjPjY14dx41ct7eT8422T09LggwmwsvNuAZzQ3erKLv+cowtKJ8Oj
6ks8rRXfE9mXKS0GJdWwSpK868bgyEzkHBhEEPCddzYe7gNfJ8Cl/pLGJ722GdyO
RAFeLbFLrDSMOU5nNsAOcC/v6wcCwLQhigW+lwzxp8tejn2HdZH46+gcikcT2QSM
qKKU0c/lpAzKaBvOMr1M2s8f5b+Gq3OAvW7izl07aWvUxI9sg2gQhzL+vnk1Z24U
j5mPJhY1xxMRRb8mcxwfrFikzGx/j9lM+M0L9TzVYxcpMlPyNQ4tOnOuzSKxiI0W
ED1Z84EHthHwyIqGoW2Rj0dPudaITmaIGLqzawitb6HoddX+rgxGQdpDr0g6NPpK
sv9L+06/UbldmQGkFXIBIkktq2kyVEPC+fnGzqs8RbMntLJrYNoRPdsYviynizaZ
mXYdGaUgAjbFbHdNbmgQP0l4gl47pwp6eCQiY3hmlHJNQuhBIEofeo+/oP338Zur
56KjXtQwg2x8BEjCmwJ5KJvMEajVUcoqF8wzTV9QY3BAN2BfuDLk4JqIpdM9C+Ri
yOoA8aIaoVg8N1EjjuQjtGXtaOZwz9Z4CzN8mUiCpTRFccPN9SXd2ckMhqi0seaK
kqTmWAsjSFQ2su67lgnLQrYSU2Yf6+8WRVNsjQiY3mIUiNNHyiz8pxqVP8BcWku3
fCUWdBGxlHMWtO+FDy53tmuk5W8SegJneOyWr7Ntz2OcpGzZuEhJDUvz/B/yucPM
LkVgzhw9D2AJrDXamosNjnCi86GKVg3BByzmp6XZMaYIoqm2r1jWfrqRwfg3k0ih
zyIKqY4L7I2dP8zXcvlLDMmCwv11cKZT1dlRyelhOrNWqXaLZ5RDl/s0Nd4FTKef
CB5ieLUM71Q9spUSsFzxb6yQsA+yiupOsu+1V9Q0WjfqXQjDjq4QLHx39qNhkEN7
FSKyDxhqNwlYm8UUN+IS5ODvJZnp53ffI22JXSg2DnyJDxY0kF+xfdsLM2pmpDWQ
77JPLtX5y6nGu8itQA2VZxpJ/5/A+0/IFrD5ZzYvUfjsI1TS/06Yn0Owb/+9KnBw
LgPh6D7bRzchSPXXkvAyItgpSoj6tRTnhsvhS/VLrGOlyrB5nC4IfDWxRTbou8ju
LoyiIgvq0+EREp5qNshTxbJPoHWGooyeUoNtcrPW9ZazvJR7GaRx7wJEQP/OWlBa
cZMMFZkB6IV+nXtfJO22CdJ4j8DuZDXnfNYJw8JSdViNCuEpMJuZ+f2gPdRZa4gV
ePUsmZiIvn9Z0i5itgp5bJ79PeY0Lo5srdNVGyPIaZaZrPAML/hoHKmNM8ZNhXFX
AwMoeKqt29UDnQzOoDCFzNs7Obf8vbstbY4X+8VLynh7CePmQiWKjz9QVX5IgRVB
bt0tDTM/HYO/QXNR16mNWLpZ4tuesKyeO8HOYqdyZEi7dY8B/JeamRxHys706svf
oQzncvbiMaIpJCM7X9NncO2yF+GCOApreBg/fA8BUG428urtifv7Vo/4b5Xqlxbh
7alR6Imn5E4xBFy0Vh1uHz8OSANARKWSsGCFFC+vb2VfuvFyPmD4gpURkSPf5yA1
ffUV5GmIdolbRgABQHWJcRep3haMT5KPb6S2YAcmk2+k3RmADjCsrvoEoIA03PjH
BDbEbXtz98UrT/ljFB77lUJV+7YG3YVE8FBnRgkq2Nd+3WkyhGOVuWGLOzhNiy6p
u8bkq6SmP3JWlv6FYUGWNNnqi0nsqUX0mk2olduONB6ac4bvKWE6viecvT1xUfXo
hl2oJfFdF9kiJOYcdsSqdD11WVgHzIvpWGMgeIC8bqKkWOaqkiort4xm2E7LCKfg
4NuEvKDAvo+FMriUsTnDpAhO5qqSok0N32lwRHgXu00Cu+33vSlObHSHrF2swcPh
9Jl7Ce2RfNsH3aSmgz79lRgh/j0YkswhrSxcs8V0WriBua63rwqgrFOrMf+G5mf2
dPoLLM5Daqlv7Sm+y6He49ZIkoTTnhoYAKb96eT/leNUarEpevpBho+RDNliqk9t
NC/1aRUA7Bg0KPyYce0XpqtvGtzmbOyLDaJziBURey78Voj6kpXSxP6ylAqsU5Lg
DHyWWC5whc/ZGQTiGkIx0tQy6o7zWE+ooNwAAiqLZUdpEkbebvirMqWpY01chvKy
ukUW9o9UAaRSZCdbk0q6xVbbuK6Xb4MLpho7vyztxlV7oCuaZTlSQsWJza7MBvhl
hAQxz/SmYbJaWLate8BjthtDtfjO3CfHDVTfTAG7hz4EZoZOs34lWpuOvjpLApM8
zQuqo7e+bW38AHzV7Cpa30U3QRvwZOQF+zYXrB1CeQn35kyWVv4Zs2pdCtbCXXWV
RgIaYGndcydJqudGG6u8MvLXwqlePDD31n/6+hBpWh+6wwo6HT8sJwQWiHKJ7RZR
sEao2lkeOrCttjI9n6RY12IldOGxFMzO6RzPy2fbD8d7qxJwF8mBPUgmlw5xWSob
u5Lw44pAAn/adIU0YxBLRQ/Fkw+57o1RrISFHcHYD1rD+9xWMU3JdzUp8zeveaLM
dRbH9fTd8Mrt1B9/lagTuiJ/A0YRFtsKe9SnWejEpMxtYcS7LRnrvgI6VBMbgtT7
ZQaAWDvsR102rgxlOFSd7bNtZZhRhwLsdSsT4nKRJYQDRk39R3x2IW7ktxTKCV1r
XDFobaokL2QtXQxTnT3PGIhZwVos1WPkypJoPPkmZsAQq9efeEzsjePpahb2mgpS
yRRGyZDJjAMbEQW9dVKy29cRmP0UZqMZ3Ai3AjLGmN5lwG1wzQzixdnSydhTy1Qk
jQ6Bp1UK5wxAClsG5ZRiCeD63Goj5yNqeBYXipUhR69FnAzxo+PyRYsTnhYYzB3l
pzSYgL6lKKsZsq6Ml3sKybzHzFJJ3JrOK/DB7u8RDiD0mfPHtbkng6fhSzbFGXvx
F0b7JbFfaNxZTMYCt4u1GL4XvAJhNu4Oucm8EfoBVCFUIEmwy/CW61ydQFdFZVFU
ZCAxikq7BO2dcg0J/C4JiGJ4WzFOejjjBg9M9YfbaOW0S4JP5LfhRNS+Cg3VKLNI
1UW4NU7XQRjazhxrXT6gVzX8zf27KynpWZF1jBRxwJSTtph/hxblDo08oFZkSTwv
onWZ62mswFHPYrG8oNtdFCNI7Ng9IachTAiDby1Bci1Gy80hano1ULycMlXMlgZW
PgSYbYJGaor86S4TC9aeqTS7XeIAI00SaaQpzHOGUblHajTI6W4gD+9b3vXofb/A
mx0l2dko820KKoyHozbN4IiVqc5qnJamdN3GhwKWVpWRdbz65L262wcQ5xEn9oMY
s6UQHTF3GO0HQtPL4DqvHmuv3NKs6r7McBJtkXN2MIlIvvnCchBAT1wcY6VTW9B1
avMGbJKXOmRJj927nxImlodAOuC9062jPLubXdtytmjB0Rjj5l8pcJRf8k9i+Lih
shlsAMXvsS0LDGsU0WEbpr3vMR4CF+8IRoikDd+GEXHfuYTkxQ0Je4dYpOtxEgJo
rrhsBxwo0hW7sWFTC8LG1vYv1ezWHBfwr57uxh4MKFhUnHYhhuB1kMFeAp4DH2DD
nCUQ0qBJuTPksJ1S2jmWcX/k8gbFVe0UsR3foNYQDVWCbafYF5GmjFagpWIAnaWx
WHN4BeWtiQAruNtf7/m3eFRUH0PYN2UKUdv0Ye7pfbmng85eUvLjP7VcWjn6exFo
MnYU8wXXgDhSQHNW7QoUEbUnya2iLTmhN3DigOkPvIERsNQdyEPGJwxYGwJT7DF+
C25Z7hsEW4BnqmuxuGwLr676ZZ75YWCqMJrctq1M49D9sF0ouPG/8LLNDqSnikGN
cPEI859XJOvv48UVPF+iFdlXgkOPTUCXvhYih/9bhRQKnqwDIPHWlvBOFI31oczU
0K4x8hDXpQ5u+wWMIKJfyNcOuzV9cJk49JVfA3MqkmVtnpPaniLifK3yhLNfEgbj
8JhCxyWVChAwCZw9BL4m13GrAIR9BcOAJqXl9NZRHgGFgkfBrA3RwTFKclFa8Z04
VlPc+QTsC+OWT6ntgx2F9B2JoH2GGYY1MIVc51GV+N0CE+SUdhsgHLqrvrxvB/57
6XD/Y6MdwMZ+Cimk4iB270KGTLusKqSQRcHBBGZ0BPBQZuM4oQPI4z2JCepPgEft
zUGxhwoRCrl8z2nw3Mf1RR41tjcKXthI7Sjg8cRcMqWT1Ob3QQ2j0Akqfpx0sgUs
GxnmpA6hIgKwcn7Jq8zeWWFe8Ur9Xb8O9em13SHUx1+KUDZ8fSwvtHBOn8Wqn/HN
1YQBC188OQKY5LCoYqNWiiBLcpnSdMr66vW91sTtoPiIRlaa+vrBZdMReCEp+djH
rMtG/5MIYb2rzPXpUkg8HBFNJ8wWiqfz1Bf1UaSb4L1SuBysS+zR80j+0L8M9Dck
4RNBpCf+Hs91D77NvkHgrRDZmkY2pn+bejKrd5XoWlnsfJ/wrkfyhCXNZ2hyvkI3
gYNJMNhp0qj/5Op8EaJzH4yKUlGmWGLVVyw9GD+bfMKQYAOb3w0LM9jT8vfteazm
KnwKuDU5iCQM8Fz6/iR0lHd4Z4DJzYyXeaOwql6xFTbzy/EGyMO7JCz4uBlFPkSM
rq1uwdOIdYSqgxGfq+KFmVFkkmdWNPXoXNxz6ONL4buZiNeeQTDyvD7P1HUP8MUC
6QSbxUj4a8XMWs6Sm1xipP6ijMC9er/qxDIhONT4hSmrP5pNz6YgkFeU7HUjVwxQ
2EV00HgfQ+PILk2t/S4dnv/gH+SUmKdzj743j6ri5ZP1C0sSnPMF4Ix7nEZXvRpt
qX3N18xZFK+mjoJGtxoZBVC7Fl4sE3crI3GZDYFaC9kjxsNgjpgid9CQ56+BkWdc
OGvLYGZFFai10ZnVxI/sp2TSk7cuGgLDgvOpbi+0Mcq599t8dgKAQ/a3hxtrCZHu
jQbGL1bE77sV30Yykx0wAsEJmvZ4wxyygZy8lUCjexHnMkelaX8aJRT44gngAUdK
hOTzwq9SrcgzKyKcwD407TZyVQV2uSK1dr8VUEGFlgYbUYF4c/Y3oI1sgnJjQdH+
O6hObo1wtYS4a+NZ39NLXIZhyxZvNmG4bteQTXGH5Fx7ugQRNRmq/mZIDYjxulnp
vNrNRFIaNuhtqbdz4FQegAR97tVTRFbDde3bKP4pGMdEay/5oObyUvmXr1jgpuDb
W47fQQXSx86enoRe7UYYTiwmr1hXbyH4vvz+43aoDcVyaFlMjXNMOq+wzchjtAmo
9E3oaL32kUt+G9njLSuwefp/4lgsHCsJrYoAdcWAgpj/hRVz+c6L+Judw0zK9u7A
YXSVKuJpIZ+fYVBK6yFhtsZMjDvpoR4B4lXaGPa4pIgaybZPjYqGXmo+9Px106lh
i++YB8CMg71QIYK8l8FehFtycgL/bfEZ8ubtUhashZWHTnIPGd163/uuRFTJTBPY
JOaW8i2uXM5N+bvmS1oKWtzyZpBaHDTx+/EQYdc5pntR8yEpK26Tn7UBJiFOLoud
ilk0P6SSC5ffVgPnvmM2bgCiMWxUnZUpz5+cBD7cyewnJwLJHr8KZcTOCTwBCp8u
EIBdPw8jdVT65cYOs6pEcuxy1L3gsw1ZVjkVqbEqbPGU9nZPMrlQiWsrLoKrxV2c
kNhDkVajW4LLJgCywllYuzhcm0T9wgizOpEccutngRQoELwjt50YmlzgaT931eC1
SSVuEL3XNjerLslNY5ZKjn2SFIGTumKOVEHdk/cX1aaSwHxcDQtjGuztJo86z+IP
lnKb+JfmCwlInRex4YJOSjgl1oosvDAX3a4v1Zadpl4gGY9hU0xB9/zvErkmLBCc
8dtOI9KnBCVuDKLf0uQ9zuhsittwkJitfCpaYY0q44M2ITcsQo4K0GcQrvwryy4k
FL/56PtO0uVaMV2gjJLbpPwQy6Yj+/PuJ78kDz6ewusp9KUfqqRYi2IbRC52DdYb
C690rO6cv9rHNRwP7E0k98Eiv4cEnKPdZqsJ97LwDBnZ6WjJIK52cFjhTENmI4bm
tMhVRoZCiJGxbkcRqdYixYdL0RF5C81m5yXqlZSvSQZh7qGVPcvx6TIEsfP7FvE7
QHifyClpcB5Pr6Y4fR0l4RU/mG2t2vFWwZRpdicsgRF3q7G6M7eRQ8C1WL8Gk5wR
exSRQw7A1cgo+edNPqSuCBeR3PjttTTc8R9hG4MOqQxcOJoVyGJIow/ZnuzsrZ0i
nJJkdyx/egnu8WYohBj/EjW6hgS4fDy0HRU01n/d+PPq9a5JBYZSETibG99g+qoT
XUxQIedDPeLT4ITB1R3x3nh6casJvHZzux6GCUS/wdYQpGq/so5sMNMcwfMzmfB7
zyv11JgQzTNG8rFjhk5N0sVNJJvwhV4DhxaG2ISzGNv7P46whWwAdF06st7B6Pfe
z1amZps+rWoBdxpPjGTseilqF9nOyPNHt6gyifiaaU0tdEGsT6KzL+il30MFiheV
68a19dE8QkDXdR5hlF5SmiI/MbNuaOEmYLFOkgx3ri2kUbMEUhjf32Y5Tmb1aZVf
f1V8rFfxWgnrm4W5fgFj91nGWRqKrEVYugPI0+Ewn0JID9y9bwsVf5weMEv9tjDk
qV9a0nA4/0IPtLFQngyympiwvT90SutyclGEHZtGuLGpsBo8taZipO8OXuPlRL9x
vxeNny+WZAZqoacZoffn4xXsbMmsNM9nRenlv0VfpX0Z50BgP0iHqmDRq+1sBwRe
p6EuX+t0EOjRhJdLQwoNYAFa0lDj53KfsouN4Qnihr+SZhNHv/qQIVzySykYVn5h
DQmz/aXrBsXfsnYjsm4nuG5H7Lr12E/KV0UlJbGUsZhrEKHQQaWBt3EOyEfGr49C
m3Upcpdj2uwj0ImXdS1hCs5ad2UTvf12ZE0SMJEybN7JMTIAy4E2LrCGmJvQ6zNz
UOK3Sj8zWhoCa1+TWqJuRouU1MCJpnAOhU52ADTsoxMLwctdWN9ucamwWj1DcGZv
E1msGuE/SRDKg/8DILxW2suaPXZvxZ8G2BQd8S2kKFwcoIm1taXZba7I2sLMTs+E
mtPzNaBKBktyAIf0s67cH5GCEmZNyC1h1LzLtWdscZPL0jk+AGtfmfPnN/BBikMx
hE7ZzFf92UQDnKBWO1XlIl5G9DYdaCROrHWCnvqRgrf/MvTJmWolmb+Lagkn7j5S
VMrsUvAgH0uZSgw2S18dfCzrE9uIBspGhXJkppLcKdeacUtz9rL538l1NFARA2Rv
I2fK2QU4/eiqIJat3kJIQZ90dcUzwqpCTdEcTKUybsWFuniIZgZTrQijBFDo7kp/
f0bP2hWpas/70uHr//3hgH7tK+7VkSEzBplG4YjnnF9/SLvdOtEwm7zQJb1EoM+n
pkk57wH56eSH8Nf6j3imcZYue5ywo8SuVEr+Dsf8Cc+V61cnv0knVR/5+Dt0MWFK
1HMRPp9hssxjm25JqOwm/yotSXw2WSOxu3b1SJZRVE93jMbXUXV82lULjKi6TpFm
8A7UBDziJ2/lBqd6j1KejXw2rewOjWdVQ/c63wUG4uP++vcWDgDprgnnvH3QqQvg
pBKUZjJTsDFhbTDdUcsi8G+i6f+QC2iXZvdmUy/ymVpaqvoPDOc9D7e2Yk1GTgSh
/Ni86PX7ih19bPAKxHqbHN91DWf6aAsNWWzfYX83bNu59gEjzcI5iuyJV1egOOr8
eN46LsJro9cBE9Pw4JMcBsRWzc5qQDykvYpjYwQFmXGMDqZkmHgmDOEJnhGf/1cq
mqvTlicCXN2es/fnN7dGR0wHRqCRgZAl6C/598dIPN5Zi5ZJc+WLfRcVfR+N3GRW
BxGYMZ1wmTuEKnp+EBQEF97RYCRbB9x9AJvQ2Nq1UG2hYekUPBC+c5FEyngizEkO
5TN0wmHavarlMVm1VlXDdsomorIz3XPXrpPnw5dnfso+5fCLf+xRw2BbXyKeLCQY
PiNvOHSuJ342NLhkSpiiY0CpeygUz4qKNmNuejzYE3txcBzhHM6N2JsouUYRaoaC
o3K4wta5ZuG5HfPyjbwnnVSKRmkmz19lKDGxlIA/MugTlxwOTRAgHPj654aqLou1
jDK/Ts6gDu/aa0IO7osl+mGwfKlGiZHb3hezda0gYrwRfo9JuxMcmEoZwwuYjeld
SgprETavRsRB+uI5iba758aCzJ3UiwPxrM81+3Qh05H2llrGxKiT2hgyMymy/Wit
7icF7DSaT1LIINz5LpW5AlIhVzyWZsWjhdHEklT1rhL1UZEt0578EPEVC6sCM13Y
i+0oRsHwzDDBQgMresiqJ4XkmZuqyyvN7Vo4fHH+EHCn37TGCI5ZVxDHSGVtLI9B
vI0ngf0XnW9gyydaKdMpmMOnAHoNZNW9b3yaFe/+3lOYFZmOUS8yLryAu8A9Zng6
A9u1FeISFuN9gRZYH2ljZohT4T7J95euqyp3BRrior3aYpKA1JF0Lw8yAUk6kCEF
dxIEKz4dSnNWxAHLaUsPygexW81JgAfZTeXgVOIpHskPbU5fiX0TL4pgjaqGCyls
kqm4I4TNs3B7ttyTuMWhQNESuAPyCWWmGDstFz14NVFrQQ9mot9HaWoYL9KT4B0T
MsuCGiaC2ktZzReYleNTVAbONhfFqQzLcRxm9L3pfN7IBEFjc0FsveRzNdlg5yfl
sBKTzf7QNOCZaEtVD/SYT8B+HyH4pyC+xQl9qF4jCoEj17pTBGDLE9+NTOmMktzW
bWKG7Ui45LgzVbaSBjIAM3O4/PC6AKCONehlj9B3V3hAhCQIapAKCoNPRXAmuPbw
wx4o+fiOGcRPYtpdeXap2moFtDZKz6Tq17Fj+BElHARGT0F1JyDT/qftzGWWXzar
ebWT0YevkCBbpVv76AQ/x7QbW/Qs144fnEUgGbLx8FGnNukupXQGvNK0N5j9N6BQ
fG2bcxi8ohCOvaFXHIOp6rM1/+3jA3CCtjfvE2U77yjtNIbf2J5Z7jwygsR6sAv/
QoJk5jwOdmogfHPTQmog3ldx7+9zCqi6F/oArGgy330NOaO3JdjRf5wUBwzZqEOb
BoNgUdoUAJ4rMOxc6k+sdgVnrfBylmXsSwRieWxRz4zl9PGhaBOnYOnvl77BuElW
OLFDb7W8N9ALgGbyJHrKN0dunB8F8UzQcI7HV6WZ7ryY98CMa8Rew4mUE8xPwbCb
9Vi9kRrt/2HHABbhFnXyECHzJD6LWT+JKskROxlp7MZDMON3GaGtSP/LB/HFK+gm
4JXIDupekdrYt2H6etzV+NiNJjCoUmLy1Q3BfX2QeZM4bwaewHIvk4w4Wdv3oG7G
A5BjIBrdLwy2X2jXKdH5/B+KBebxcJz1Ye+ccao0KXBpr/3ikTuH0VIW+tmbezaN
kOsChfeofGy7pYnBvhI73ijYcmYKKTIotVCXm4Y6JPr8cLGc/yARrBwJ1IibkTWS
VNBYmE2rKyNwLksXqzQ5asSHBSmItfIpqNq1MoYF5lsILySAV1zyR1PkQa4/5JLy
YEzI0XwcEAhACmnULMgP9+IpMmL2wFTjm0TcediYjUnHIhRdqtjl1YXPdtA5DuwP
co1KMXCPnVv40BUMWXPhzO3UDO5jcvXsT2B3IulVquEdBCfCoVM0W/SEwfiyeVnK
xKbptH5qGIwHSsaikRMccdxbLXpoMCobSlhxfSXAXv8S8FZ7gjJveYEA7w9GLhj0
TVxZsYvyH0E8sNNJ1KkfpAbfiJ+NF9rNe4uqkzvFXl6FRzDyj1asmRRgVXQ4V+W5
AhTyxE4AGQj++HYQ5YRofINj25xX8nFZShUWul4e6ANOLIfNkHMDGqtGfCJxVrfW
iFREgK8Xgkl6TUPf9ovlmDp36cLeCVPUxdcqk5fEyR8IMUY0DZ2bPNxRN2Y4BWdv
mzxkv2MrI46RY+lW3ExPlzkKZkAu452pNHzWUi3zrIwHn8vvvaiTQUjf2t5gZS6o
yUmvXgY1LREtVpTFdB4TmWvr9hLyL6A6xjat34GXYligG0fiQMjoUS0+zmeQzVd4
sTKk2xj1ozu0ptQZslTtejMPEBb9vOJLun8h4DnburMaTN3xPusGIj6kqz/aRuJl
g5XH/zCsb4bIrTjxGf/fHDlftkMyMBjL0ahy5QmyTejUPzp/a5eCkuEwF5XpRCxR
5qqYgd1Rvuu7lmBUDs6oY8ftELdWDIEGFOnab30tLj02qkZdb7hvEp05MqObxn8J
a1OmS1Q2O1eW6ZyQSqVW8EVzSzpoOYRD8DCCSll1Xom/lsQcftcQjcBiPxHG/L9i
s945qxQhDpCVVv3I7qaguTCjg4XoEnJ94O+xTwIYYQsF0xavh72pR0WqopLKnjn6
ymSl/hiPduCZFZR8CYiUoV/gRSlI2NO64FwTiYo2fVenrrB1toyaa2fNdoGD0WrB
dLgblajCZNx9t8ZUf7/w8cOLdAhfFSuMEkg/4OeBd1g9s/1gKBtqFyTr5JUdGWWI
J0eREpIosglJY5OeKihoPxRbn//v3m8htWsufVmX0hYQjAlPzPV2sBzI58CpntqC
eHLvFDauPGta+NYb90LPoPlTwhvWR1ey3jc3c2LDQH83qP1EPWG3EGck6PFl1xEK
owczKGKUSRTyNmum/dLHaDbUXDvo8NZAciDvC4qZRyTMwb8vcUNdnSFrsomz5ICm
Knk3s2L7VxJ5UReyoCALAXJNVsgJm2j1GAPzU1K3YALyzwNDzHxTXWytVaIvqLyx
EX9odi9d3NUVwvf0RFZcPwDPKbAVUSjkVWYl1m1b1ku2ymD1FbSuBgQWGEY3eycX
+Ct6HGLTzMRU70Nkff3Ft31rUDh7rlBk4EndRTVbFKgwAT5N9SOX1HiMQ5aHIS5M
zlNXSnr/+eHSyIiZ+E8wCs96mAkE2pAXl472eT0zkExB16JPayB/G3arcfnB2rXX
TzynyfTJZDML6NPnYs2lE7hU08YX73MZqhDzz/ck4L6YCwQFiJs6fRYacD5LenJ0
UPidbX2k+RTSEBB2FuImsU/sUrfX1RaQUbTHuGCYq5zDipotEfx7HscNBfasCkoj
MEZ+60g8ZCtz26rsPVgusfYsfiSFjYRyBnOHeAN4O9h0TVZu+07tAzVIYgY+/AZC
hos9ndO9RyreMU+7q3M4EXDZJlP7R+Q26RmhFnZDOWfccr15HybtG2FHVorux6mp
jOxuWcG4InPnezuNEnnopliuAPEYtCHYM98z+2+n1/cHiLvnyNxqJ/OhT063b9oY
4emrAKE4/DUCi7e4XDva+8rsagxdTze5RXtAGDS5lt9xQVYj2BBeZYhYyexFBWPP
ri5Q+ebaYmuelQmy6y1lv15w6/paA7duQNbjpwjq7cKWH38cEA5IM2nQOaAMBbLD
GsXXMe6IOI64s9BHPPoSwlcMcYZuDg1/7J+LJTbkHDd/X5H23Kc5/b5ugUoLikuF
v3cqDPo7vPDUIk1cqqoBK8VyMPBm54LkQA0vD1B+qC3kqjaUsr5A/6BkEBbQs1wE
B7HGJgt9Na1rA28JADYwWUDXRjzU7+wSsdZkNXScbiTtbBSjGA6rlCAar8S7dBLE
WcXfT4xyg5jzs4Xz+qXxUWYfV4wxxoVGPPFmJ2e5Frwd0L2nho7umqBDIy2qtHLU
E5R3YZogAlFLmjRFwDZmPL3acoHjQqgB7t3FJ0Rycyel7N8c9gAY1To/AXWk0jl+
8z28bpQThQ+ZpEf5UmjYew0ezR001SK8Ls7w7+lhp7IEZXsefZ61kPgTNbqn5i+4
57wKL9NN9BQ+EqOe1nIlgjgxJng+T/4vY/9p3i+KZhQbXy0id7aDhsQ/c1dfu5RW
k4SPVQA8+VYVmqipGXDvtlbWzvcuabBB3puevXX3iBkgsWxeL8jym8HGLoAHxK0r
mgS/VtAXSSG/xFTN8nPUN1ec6hztWQ7vJwlxm2neB93USpmHrWfTQi+piUa40kGL
qQgAGmyO6mtmTdpOE04A1SlA87HRNJrrcsy6oXc8GQkhtELesJOHmtGwfgtPAQ0h
Zjc3UvoLhQHGVLLXzj1Hvn+EpcqywY6C6gnueG4GVNFNMfyb6KkghGmjt16CTUEH
nnRl0frw+JNEiUL+rnMAViZIMw5ze5FlXh5GRMzTr9HPjQlmjjK+CpC/DMkod9sI
pYVj4GXAB2fDIbVQyFA0Szsb0SorJSVwPRRX2FApk1ulWCXQgvXHoD2lWKqUvsPY
wkjnwOkWIcumR/sSFeb2hUg88/uuXz1xG12KsS8ZTfR/XG5F92dRagbxBmY224iM
4KnzGLuPsViijXSceGIUkvXDEkgaEWRM8ASNEcGJ+3O/hAT8LBPRs/J0OUFsA7ek
S4vZrAdy0Oz1ixgrHDSLlk3Wia89cQ4HY1/GUwxf6N4M3MBwzJJ+e/59AXRJ87iN
/VL1445jEXeWWKz7F6W+SHT7a48jBIadF0Ksd0foIE8p051Xt4HOxB9B4GRk6Ggf
dFha3vyfeMpS3WQ/FLbxHmZuAt51WRns/I16TXnk9kLop3RL4XQbxJwzIhJeeFJx
TjdEgR5NAr41VlRL5I1U06SYJ9wz7Kx20DmaLw1fIXC6DjjD/LFNECI/5Z0izH+G
UHdKPt8yiopiWQwNPKYRSDI+O+U967wGvvx/7BIxLqoJYujbMNM4Vebg1Jbn2REd
jwwaDrBWhMI7SP1/Lw+jviROrJq4l7GL+4sfTwT8MbM3047hRF62TwMp7nQCKeUM
p2/AQ7KHzamdRu8RB4Lu6f47WjcqGn/aN8kap31azFvYahJK2u3vVsFmKCE7VTAT
QTuFbBOwwhOXaZMAJTLAkBB1vaU2mBAnAM68HXt3T5hn74kBjnk+3cGsNpN3ZGXw
Lw5BVwfL0dAZGjhePFvUHqA2CKMM4APPEonaDU3zlnYiBOYCyfFLxOFiw3bbaAww
DARxvaGbrogBKO/vVE9QBTdyMBWOXarXFw/ULSJ20CbpFNNuh2iA2kJsgqd7wyNb
vN5LLgeL0pKrRmMtPz/bpGPSNvrRSTJN4Ii/3ZLaPgA8jksksXRjPGhTABizJshg
UEhUE+U1ZctQ6HxQ34gpkR/V4gdSq9Wgca3RHtzcoAMnTQGJGf8l5vihW3c3prsO
GejSK3silvSnjJWCqq3y1MLyn+RG/JEV8heHSUu6s2oBOiidHAmww8SiUG7yApuY
x+AXrXfNwcGt+Tdj/rCJ9NCkf5FcfQlR7wzVk1XLF1SFB5BwLtxElRUtWaKjD9Q4
xhNdSA+qNQ1bZg3ETdi8Ggk4F8j7nEskQ1DOWKHKReYUIlEO2KG/t485BMNnkbBr
O5ky1EAkhWTOXPHiMm0glUeO5kJL6lh77YiccRxdkphuA11J5o4Cl0+kIqfBgiKg
rcg6AWWdvNnHgo2Frwb7ejQ8NBI1qVx3Aawmbs0/oJ4KO1n43md+A3Cb8EbuTAfW
weBW5LympfWU7f1Fc9aBL0L/NlCQUc3RDPGTmrlmdVmaN2UaCbBpWJ6ZvYAZIlsf
dKcNHk7W5oqSXJWYqgTVUZUK+EizseQlOWwJznYUmgCHTyhFuBgOyvzc65m062gT
2ajakvMVa2BJkGBTOdc4Yg95ChoLWXon7kaczspklb9Qpzn8Vjp8g8N+vWHPgK0R
RKEj7YpRQq/ap6np4VZCFmpPqO2+gXYP4WayCGsT8NEPdiC+bdE8aBvGbGCE4b13
UhPT9QsJeMsBqHU34JT8ByfMuLx4U3BirTbAbmzOCVarS/2Zx3PfSDZP5IIOpbpV
T9yywDnZI9ScUKPtLupws/ZDJznuRxdsL29iqh/P9hwjvGKMxbus/sabf+NEUqJ4
yd6o11Z1BAhwynVXcgCSJNl2UJWMDA+h5iVAbhU2WvMiqT+L+NfNs1NUBoDjtYYq
df57toeXAmwcwRGG1LtUTUqvQ8r3fvbYshrAZ+L0Dg4NDl9SQSh1rUXkgXSQuNeK
/jX8Srn49TcE0ReWlMPz/dyAneJvNAyYryDMwoIw/mbguSjos2W472fFpTjlt6um
OaMaCpGc2Fv0BIj45/lW0mZOKNhv1MDfVPsiuX7VThykENetIBY/lDUubmzcCo84
8GupmkaoSsNN8/Ps16xioZFiCXgNb9/Dpo5RUcdvIEfF8yV3oCIkuWwnqKAzkvOb
PxoEdCro2gVfPdwh+eHCTkHGGi3HkxgjID3S06MtI1HeIFSCkKjvD4N/4yGqSL15
gSlkbjKaCRKWEJa/28ldjCSnmsVaOvZFBSxNYc3OL/F9+dg9TrVZxGL6wCnlPWre
CTEO6tnZUnYpLcQQd2vWDNPD1FCjk1x84pXa4Jh1OrK9RPzpAIovmZ3SkTCadAFu
z2/1tVDIbh6Sw9QVoXfGwxnkGTS3BVZfuD+IK1IkRk1ye/mbzkBciKA2c+XG7X3I
mzLzPbugnYM4nFqP/kDDVtWWgXCTrJBXFO8ONdHWE09yjttvDFZfTHJdTNgB09P5
87Y0VQw1e/aQ/NczH8WF0dUJzInkBRMrmy5+Pq29ng+9kiwG+gK8WEwAoJnmuqBu
8PuMNH0yICFX+lJGGZlwYWdlkj6w6oOXuHGzpLfYWY/Yz5rvVc8Tt+SX9kTwwmHX
pZeBxm8aglTn8XgSAhlcn8IVYqZSkn9pqdH9uBV8slc56huw3Uvjp98uFJogWNaP
Wkm/YFOrV37miMHs0QGhRFWWJk48QXDE0v/KFSSpqR6lTp6dQYwtmcb1VGSvBO7W
m94mNA66ZjT6dWu6gvGxBX0bC7RlEvxmC+V4+zziPgHHUxKYFrU9DAg8mlytNUu4
LoU7YdSbVaLmH4n2aCEptg7S207GdbVasZ34p1za2MSDsTkMX7eNikp7ZRkPUNWg
StDHip36LJVVJsxtnZygfmab8T8vhFoJRB85u7kGXk8o3/07sF1elldJ4xqtqKel
pYQl/4dAkPG9zLHShLBM1PFond0r0WHYkdKSR5cH76Na5zrIpuJwMID9ouTUh5Hw
6Dz6bTeoiHRCpHqMA0LYpjNQSi+xT0420nRiVefBSq1nYN/vQXCvHilXMqPrq6W6
hzP5bGhmlCgqhq7Jqhm6jYMDlgHy7K3lXWZF+BKwJieIGnJxL4cTw4oBXk6XgVe1
Uxchp5m7W8nCUH/ligyCFs12BUbWn8cWCnxSXdpqFKk0yYRbzLk2+c91z0qs0RDC
hPwFcsap5QAlDnKBJrxMb8sggp7WBKDh+89CojDhSzsmwBXF5/O1tmH4/gjJntGG
N6EPMG1Ywqgu8LI+1kzmvc/eqbAkOXrFnKGUwUi0I8pyNKN0p3o8MAuFoLWu/YRf
v7T2sB6tuhOuv8Zowos1VZaV/NnhrLcQuWdoqP+2Z+TbBRmcq/+7U/Bpu+WVVXJD
dqm0IL4B7pieuvgIFYsxQOLl64mQg6ATUMWRLZ3S8SubmpdxhK8YtXjUh/vnF/bh
INeosjN3LC59Glad/FbSfyqnR2LAQWLTvwfjF/0pJHOlPjiJLq3us7Baul/VgwLO
KrTe8Zv0IQrbDYGaEZTI2LxsibkiDvly1PaXEYKVrMnhEaoF/F5jU65xGjqMQpNe
amiBdvZHaoHf0FdF6IVLg+kmXqtr4PAUsW9ckDFQIA+ZDaMjPOQD/JMRwi9Us0O5
UeqjDaZvrSxUkKlIWWTpEx81AbaDfUPDpM5HVpqLvG+FRMaDwSgHH6t1qVCMqD8c
+BJtXmBJU4B98EuQv4dwgtbq4Qz9NyAnAHse0/xS+ariDyPtaO808bQF0wZTgJnU
dii32Q8PXc2kdirrp2VTuLlnRWgtgvLEoQPvb+9u2njRu70rFBSHbGBFn3eZtY3Z
2u7nlNvdHDkE7cKGwsofAERsoxv00bCk13fMNYGfTFfQqtnKWOxMeN98Vylgu1dd
8utIk9nH+rxqLyJPaC+y4fGOk7lI6l/H0sRB7/eVt8OQg2zJc6JohBRcHjykchB/
0VGpn2TNE06fZcxzDTFJKY1FnkOrz2zHB8Fs8U5xb90YWpnOVLos96AQappCu4nL
6TnXnHjrARf4m4RmNcK1srqN9oo6jxFzOpAgc8qwDEIQ3WGlCcWf8pXewlbZtB39
kVWAVKRmNymjqpNtU4tpW/c6rZztEvqotydm08/QLEePhQND1rAvq3QF9iCzIoLV
Fl2I1YgxW1bHHjBjFjdp048K51Zf2l1/jid75pZPi8omWMFIIMFBYMcDp6I31nj5
8B1JVxskx+2uIo4QDwHrLYWr5teQu/wrrYLUUdEJe0A8brf2x9ekt9X21RC+/+wL
u8+inx1y8LYa+DG7n/AtMUneNvDfO9/LlthjDiAJ2U6uoftxmuJgbaYkzxINWtMD
iYtPEuhV93wFxDeMrI+FeXou5CdXktD2+SL9HGKvpDKRZeuarKOWiuEtycuUhws9
JQqCluYEvspwgwncdQCNlf/0meOQUzVE6at+lYa/Wnpr+M+s1Y6SIee9HrlYJ/Tu
XeT/ZAV1X7Q/6M1Y0HWu53iVjVoRkbZ8dsGExx8NWKp0/BCz2BdH3uQoJ/UrnQm7
HG8217/EkRVu8ut7L0hp8mMoe4BA7JUjk2ZZ2QeHm6YMWtfFWoYtplJ7uPZCJmbh
BhulckJqEZDFDu7d4Y21fRtgrVBhJARZet9xSakuG11eEJhSkf35pbGg+TdkCru4
C5VfMyRofRndQCG4VmriyZbakyD12VlE0uLeYPj6zifehEPQWUSr9ZzF8laYLCA4
VWCJPbthusIDycYo6FY6mAd4wx3jGUSL3RFVb4MCfvoNrvxgOaFZBUDqRufEcdqJ
rtiwVk+lNOizGjIYFwQZTSPIxMbuPEAup3FgdOddY1IGxlvK0HM+K7heF22Reioa
WkEoUyAUeeGMQkWjywVYKX4lmMJ4F8X7OYuQwHdveeuVWj9FIomPH/V55iYP4fgo
ojTtRQiP7a9UwYmqkA72wJSvmTQkJ8ub88nuzn4mVqQ55Wquz5KBKgCDX6zZvUKC
jZEHRSkHvqoNnt3iNoiW7MEWavGwJQRvnnfGRyIppcTPt/a9cLCpGU4vXU6XwvQP
bq0uJpGV5OBiZ46ecXAfisTc9rFwtRiEJsPU43Ff+o0aOPU667covkxyZwgChhl+
S7oGIXTjgHpgLbJ219Iet9N42SWNR4x3tZrWcT/sJgRj0pTYs7Yo2row4rDwu8xh
jYHDK0xu37cDhujsQNfiUFMKKg+Pbr6lwsdVkEDfK4tt0MKQfx2wHVCf9/D/aHjI
3/Xa9fEyOjFRNIR8sVVhin68EyrrMHC0uawtbnZWSDT7CPhTzjCJf6GeeQzfpiPW
btKWEi/0p2EzFTnqOSvDnALPUSnixMBRpUkYCznkA5GHhHEWJH4TopNu/NCtetSg
bwjhSIjREUILBaTaTqRK54zi+KUZpcBHfh1qYquEXc1wA8czfu3oMrtScydysJJw
AUSB6qtPgqlBCkm8jYt2fRSDQjsQAol/qOoJlL5Wjse/CqHqfBwl6bozmJHRIzBf
jRFBBNsJAlPRw/Fxx0rhfT3TYi5qroDJ+CyEMUiSrSltIROORlLVT0w4FCRhQtnE
E9eWRWvIw0Z9KzvGtx3QzlNfn7Py2pyFUXCV9lIrCTHO9SFXCeh0CGaeel1nlT5B
6T8rUTDIuLizXjv92uPnGX+b6osIgM+bL+BV7EWrXAVq3+ePkDsc8m3lw+Hd0T1m
tW4Bl5rryjbmkKyo6xNbRuEQqKVZmP6gRuD1EJs+mAmspq+3EPW5PowABCVOrYjn
eP39L71bRnYkPI67W/53m7xEHxPVFYmqwndRnvWrIQhkRhEAinRT9YUPT2bGz9m8
dLzvFcbLaicOETcxZ4BMXZI0/ogGMLf3QO+6FuF8jK23JW42vhACc8PRoQ2W3Z3U
TgaAyeAzP/Qk9nwZ2WQkOcRwkf4D+6d0ug0YOpcTiQbI/qRf6A5WcUL4LtQ2JuoC
OCW4gcfVYeZE9gCUaeO6qFIyHBZQjWmgTp8duCzjLknZ4LPGDb8zDWK3I5dtf5Rf
YuJuGz3F0EtCbP35JyaNbQ4+F4QDY4h+viEchwCBIyO5U3DmvQpGLLK20WYwHc9Z
R713thwX8YS4xmGriaSAwwXJNbx2PLdnmUnUc0PJX9hQu9/eaZsfF1ag1scq5iN8
+xjay+yGgRvbtFBr4kc5rnox1W/hS+jMs1rZLlKfu8eCIoy+I5na1h848ulAcZjb
lu3oHGpED3RHYvTmYnFND8S2vfOesYDkFmMxC45B7mpcAJoJCuCQY+dz3lpJNhTy
KPPuXA5EnxnLH49KhTfjxCxLhQhgiJAZkla2JYRojE/OYd3GHskRiAadnMEuwsna
8I8KM1k/KHJ4gkxhhpfu7YUMA65xH+GdowkTpY54Lo7FZ69f8K5bWYMbiaihdzub
K4rXu/1c6RSFgMIBk+T2Gcub38yR0ia3Ob0vZUtPyZxNjnf1mIlSmtSwUfG0eiuZ
JcatvL62sUVPXKSppoRn9tlnie7Pp6zuhSLQOGRqafM7/D3DhZnB6dWw5shwYRXm
xQe32X0Hj6JPBCiSMtKrj2K57/OQOAQ0/G0rsoyc1nBu+HbtlfuTLxQNQ3uyhaB+
7GMBDt3tsWWaS+LNYg5A8GdIRTFv1GaayJiOVk8MUN1g34+yMtR7p8q6LS63OavP
bQ3KvV0AiQ/BGfARz21lWqZ08G0Y54UQNp7wZQRUtMxuQ+AdGGKonbZJdxUBr1MJ
fnkmKpuhSOMMD4Vh+/EEyzuQrWCqi10iBLplSc3/GXPvCt6Q1jDdv/pvfYjNTI/E
RvXX6fj51M8MwiNlg/Kj0U+PE4qfx0Kl+tGYE0hbICRHBOnPU0i9hBAF3rEaMidm
LxcysccIQOb6kY+BT+KsAde7hANSZ1oWtzFr96FPTwI15321UVocxOI7HRvvfBfm
4gSqHz0tk9xJ9gHSOjUof4bwFAy9E4F0Kshu6M6e+s2wSdKL3BNFXG2L7zDMFtLi
wEC2iW3g/yU5DiJFIh60/7+Sf2DLQoZiF+eJfXBuV7c7dfqiL9chqBO+Fw3qP85l
pdSb+RlGAa3r+KIaTAC9WTtwh8Ey0I9xT3ecgZ22iGUqODU06LKbl2Hz3JsiXrZC
vH2c/CM9ODEB8w10eTXL0tOljJfsv6cNOiIYecSedMtonU/aWvru4cgx+D9EQ+pe
IfeGN5fywmqN6/miVZ3CsHbL4csGa3fi2wlsiTQJRHLlF8Q6P/b2PXQLvHm0GfB/
oT1nvJPj4X6gx2U2Fmjp4m7CjQVxeQSom+miP0EZJ24sdPpNRRBpyYeLnWYN1hIj
tnjPWEBTnxlvZxhsP0F2S3UQZMz73bjPO0iomB2SIhZIJtSinmrbybAuYubqxDWa
CnvWhH7d+WwWsvKAUy4hQpVC1J4RQAclnWTOoflr4DPeT8CD6ZDpPPWzW0rdbSr/
mOBmL2by55OYuXeEKJ0g+u86CkSx9FabsDtLo5FMQ8EnO/ETlZNWZkuNS3RbVluP
lAkd7ZG+dR9k/adiLrl9K5venxpQQ9C74MbEMWuubFNPnwEnfTdOFRGpRlA+tJ54
LRX+h5DD9GMqXwT5VHSTr7AWpoayJbOTlCmUW0rSJRW2M7cNFj01VMkJFFMF7lfz
DjFgYynqN6LP72hx8r6Qz1ulNh9e8VM0EbOkDESLVI9/khPZ41P388FX2weiAJ9F
sSjgvMXWxewCKEJ2WzYItct7jQPZOAO4uwSupeepA7P3GlQUuYCqIszO5SwWFhPX
WRR6hLpu8It8wGuyX1f3TNVFtI716zWkgFOqLbiJfOl+HtDeswBB06HsJGe9iHCO
Zjx60bwhVGgXOClsXw+zXFLGJmc+3wAmkeUyHv8rA4E76Ph1l9BM0EU+I0vtuQNv
Ys7gAjknSZeO7XnjB+rzmS44kbsA1XAc7xZfMn6WevgVxADMNpwnGXuiz3Jr7Hal
U71F2XbST2VWHjK5OGuCqp8Gq18oAIEPshuQOGEBePHm1U1pwoUNFoWXhQFJrs5c
OXXsEjoDD/kDem7EHAWuBd3gIAFmFcNvyT9Gnwb0rJarkhly+HnbRbZenWwmxM6u
/FmvXATD85+NG99uskgKtH5Xqh7DXitdcutUTQ2gLvXENvdBY9adDMxfTcofpwBT
uSOvKiXedKf5BPEJE15OmgJQcmbBDR44Tw8H3psh/FaBlmlU7xryBlJvumKaO/Dv
EUR12gOwUd2yPf2Gcsk5m1Ox44KZywGR3ysSqfSHYQJz5tORpj6XvcNE5OOhdPpr
qhtjt4/MCpqSXKshu1qXFUudnPsGYBcvM/N50WE2BGB5vPiyJI6Ki/0Po4K5dczf
Cg237YQPSQI6pk4QZk57bA2YB0Dxy7GFXNB6VQEQYjnwpRRzGkePEZ8fy2oKUVb8
2XXeyr8ph6p7AJDArz6iNVbmCAQpU5n/A5NGAGy7JxC4Jr3vDzX0R3pevX3v2O1y
EM55A2IX+Y6TR2QuanjCERKBlnRAPvmLC1PUkDDcbqgQPUxgY/9P8+m/+wlCAjmM
JozzJ1Z0Ppbyh7w9cH4OwBlIl6uB8vEBurCjLU/A8sskJbqHD8kZlsb1FcVEd1Ci
HpAhK4iuV84tVjU6qQnqW3yauORgBuM4wsjZD7MTxgwhDa1LqZ34CdN1p/Wx9ncD
b9vaMacjG79VUTgq5pZMhbgvA7vktSV1LzxVR9DgZFQN99jBLtMhjV83xIuXmNok
7Qua09zL3vRRXLWWPauaLWKjps0od+PTJeABlHW7sxVc/vSzTTSzR78ud5/Lwbks
0j4xEYAhE3lHynIS8r5GRkL2hUbMNBz2Rs6l0NcDE+6ikZSl2HEmmv/ReKS8dqf+
O3iQM1/KXsveg+JT+13/vyU7JLUY6LCtTc3+W40Z2i4tRfkMHMOewuCSMjpwsNSu
v1tQyfG/t5q5WfkLURNwoHk1JraGLfYwhcKxQlAA92HmV9rzvBABsOmu+NlQl4cx
+SsXM9tT+BiR4fR3sFRh3SArEjHKpDqrAgiTxeAmKc6ot+FZxXIchMA47glfMlH4
6nZfGqa8wC5wtETzIu/Du9pJQp/UifjAdO/HMTmTrnpGNUYDdBLTxIjAKNe8sacn
sWB8hKjW7inHAsTCspo7p2lCgdJKKILis1eAGaK6tzkAs7kstxkY+Fe1gJPMifEr
g1cUU41Ra9SUxvy+/NNnuu2rXBWELT7y9rrgZaa5udWlj1zWSlzSG6u6oDnJu9d4
YDy7f0y3wxLLsc6lkaimFWLe0X8qsEUtAKXevGhzzdoXnebH6HP7k38nMn3moY8R
6LYpcQ4YkxC1GvAdJAJ2HJpG01/O7x/NbdxxNdqyj0TQZfvdtvTtfDR8UBRx6CUg
N585Tw6MSM8t7sNqk8s1flLPZvNQNLNTtquqiyG1jqWC3E5KAekAt944PM6a7vqi
ft9nijFixJfwq3bMgv59AEqkCzUXG9BTYkwlkOhC7vZ7BlhWWMP/nlKivMH5nMIr
onWw4kUbQOx1P+axXuWDdSIl9jOn51niLP/YeF7rsxWECx9UcT6CjcDBDAiHJ1+h
qVOikcP6udDJ0DdrcjziSPLgkqkN2+ARzw7NX8HzSCBcMR5KMx7bKr8ldAOJerV6
z79rxVdE7/J0CTYoQ9Mio1bvg77hSMyJmfHHXzy/NchVzHYHLNz/MOmNHh0fDyE4
ww7w5SjikMNOJUJ+GQ8xZW9vO7Yi/tSSKRXcACHsq7mq/3rj6xFJDkKOX1jn+QiJ
lnijUSB/ac89OkxsoLacJSlCG5PtqdRkkedZqFO0n4rpA9eLFWDlqDg89NnJI24f
FCUWE4jyGW+b34PN//j/R94KHkXN4gbajzW08GoMUA2hZN1ef9uZGXKQ/QMQgl2o
A+sgW/ASXhe3cYWElsiTiCLnZn8ZVsRTz75TMeFPjbrX3MK6JFnfVP8nveVu7uEY
luAVB8y6lmyEc6rORhw5en/IAecUsOe+NMDP4tqNA/YnIRdQ5ubQMIAQvzyLa+a1
l/d1ANAA5qx45pOBbxmrj743fg3bE10yZNVTau8dU1VgKJQGk8u7tldfPD74xVCQ
CZnVFlsMZ1oi/gMfRKoMjlFsyawIz72AAmtTnNhNb+rOOAiwu8LY55gntDwEcun2
tSrteZAS2+qmdWTtfARjVfelL3U0o1fgRWapBf0VtNJXWsIYpVI4pjvGp9Qss1ld
IJKUagtgM/F9kBheB+fZYHflfIpbSje8C9Hs5t9tylXS5jSwaagQVkSBO+ggAv5/
Ame0PtiZ0QCJgAPRbuAqdbac82yv+IPvx7IPQqCvdTm6wEAYl6D42jbiyQ9GTAX9
XjSwi0YBlLzXbWLV2mZtXmG1NHtIsVNNEOUB8aXymZnf8kE+EVSdYyarBVLm9HKz
lZDmu/k+xVRmGi1VC0Nw0WgK6wGv3TNytRK7xfMN21wkinM5x3oUJWtV4pp7izMG
Nwn0shU7hlzu+vEiS2qiqVpJEof5vT0pPFhF3GmqlvgjVgsE5mZS1EYvjeARYrjR
+D1shSsGE6U0fOu/DiM+NwBII7vilS2YP27P14iiZGtHtoRZFnGszkpwOfQB4VQ+
O6McN3gJXJlQ99R+QQWOSooG/mmRz0YP2ixBRj6zX8y9wzHg2bpYJJqesqPY6eDb
i7weZA26vjv21ZQ/ivQa1iNbW2W+3ZQTrkleg8NnbW01lpdiMiK3ii0wrjsP4aEu
zjpdveNQvRq4ThTHJpADyDq/OQZh9GoZXlq0SaqmuRX7twB/IZVtfwdUhrotJDcM
0KVrTntzJh+nilqRcG2RgLm1nbHqdnM8SsOletqR2T7kUyvMvQZOOWaBEe6gajrU
PlG6Sg7LOq+dmZlMHzWVwWh2OLRc49x0MAWVVPBrpiVjvsTMuDeH020L5wdMJKoc
OMU/RC7OmSeDZXU/bY1rtvW5lYVdu2uwDW9FLldicZWLT5SOrgGw4IhwK96EJIB+
2I2lTCse8WhRk80539wjsFbzTSH6XrB/MVU6c0AG+81NGrtQLHEeZ5s2nc5A8E7X
+NryZlPD00qyVhul2mfj1XHPubImnMwddLXXtlAIFyW0SFwSxqFitgnJU0ELFUbA
nlSs6+vS25KesTE208geA4F6p6yuk4ALgJ6Us8p8hSeOcKNU1mBZbMeI3ITD638E
vbCRZ54y4pBOJPNOjwYDiDwjZCKmZhlL9qvZwGUo+3kmQpy/ZVjPUPCr2lRwj42f
KzclQ4ELTbpTSijjtkeUq4GHb+Bph/Jy8xWCiminPM9bY/LlvyxZcqFmYOwBHH0R
fC+IAPobMJCb39uxqxicWhRnw0I4bVZnzEKTz7/QeKGKLGN0HFXzUFd87jJT04B5
PIP3yu7rx4s8ovK8vnCn/oodNBwxJoOBt8BhOSHx5F7NBxLlY5OVrGUF1DwlD+d+
AnRMFphIGNOUwLTnUVHzejEZsc5PDGsPBJdTe5GzV6RRtQD91OMHRvSFZheU/Ftj
ZaaQguMPVVFatpy+t8sdTg1KeMiYc9YofltmMt5O4KiaZIQUM7sezmRZaOYaXR3y
ELIEBkQfNFn8+pidAdQeYMvSL+KFafoBim2peN9y3qtxQSU9blJa84HEXYsMeWrA
4i/CxVbs+YNpVERXtmuxtjVNcidFtwELXxUucmA7/iXG5e5Tu8/k46rhFqFCTmlM
tRUstuO2ujkJzP2eJEunb4zSuGIx0JMB8HTzVtm1CERQpUBdWlp6iX3PkoU0jMkC
jATTlGp32TLDAji2KLh83OHPveT8cV0RKnVz5buXdPaPU9APG3bfq1bHJpn61DsE
WHwgvCv2fWa6jQwaN+pgPOwyEBu5K12GPD7joI3zjkoNr4Rt7f1QCbwME6akdoUA
d7504Usb3MHcTWPN42PCb9rFLW1WaMww/ecNFbVlksT7XUX2XFhrfWgzMXzMIe8q
011IH+kwrSVEe2LGHNFDWfLzDmExALNsfq7+ibn69kTBYsuWtnGSevxny7/3fHzT
Nrw2jDiFEM5GejGPAFI6+TYZIe6bfJhsyg/6q5j02b8gCezdPPXkkbULuKzmh0/4
xZfRk8KQsha4QYmouAg0t5aOIRFxIIf45s2xMVIteBWmV8b/EG7qyHADFNCkTsKl
DNFb6nRWnGySMhYJC0ILT4RB6uMo9TH7ZcsaeCDuVNTPvHnbFuBrpDDdS5mkJQX+
TsJcV17aeab3elN3CqdZj9q+1/8FSau3g1KBtt54PMXD5xv8ZNZMy1WGlR7beK76
HAXx3rrvSre9FL9rie/qFta2VI5a1LXT2n+Dt6trxqPOLysryIT5KVKBtZ8jwnW1
YTu2OOwafD0milVRPx2BBGFWl5QF5k7vHpoNd1T/m4MiKx2MSiwuTMCNZDvyauig
vJcBKmPNOk9iO3msCUQpMvhWA/3tw7DXBuzjlixXt03uHGtj7EfobmjZ0+gS8xdG
+CoLboGM8WHtVc417vx5AEQ++mmcALGS6HVBbgg4X2u5JjKc5vsFHERftLjaBSDM
WP55sF0qifIouGDVlR93JB4wqLgdVIPdtZwj1l+YDKtodqV6WZQAjihNbtitfwMt
V47IM/B5YoYxBa17PYKxrEByzDAou0smWvPss07hkZTNEwX0GfrGemWq9IonaRXU
L7zoG0Ufj/zPQjcbCGI4x9vHnrdVzDebdYRfw0yCSQmgwlCGnFe2kauhpfZ54gtM
3yKpAuP4j2Vosa4CMLgiShEmg6hPj/sV3urvR7KL4dQgFtrdZ+ZQs3a8rV8qSH/x
fm4fQNWVs0A31Flan5eaeSgEjfQ7mTy7CCtHJYY45zqnhqzreYT+kkRB+KnDGlto
HNVbhz3JvePHbDY1G5XvXa/99MBCxWXwvl/SlePibItW8XCJavOmM358XBEMJwhu
/vnXDaXoCSufJN7Ro9+apdvMpi+KSNkirktEPyOpjkZNFGltmRkzBgIEyTGiO86c
BXfKFQVGr4w71JdQChb68Un6oDoytB4ojGvVmoGAAHprSBG/R0M8SI5jWlSAzSJ+
8SjPjEekHg/0k5wKx0V/7IdR9xxBNgYG4GnSkkbThywGdC5UWZyNcxf1e1IhO+cC
TrB4mSBWngys5+hpxY0q9THO1iPEJ/gukMjDW/p+DGS2Qhl2++7BsAH13uiG9Ux3
z0cN0TBypCoAOsoaFIIgT2bJwKiGgwjSEQAAvEXwdVIhWy3JooFHiv01W9BJtszM
JJayZeRONHjtYiHWL/hdeCmtK55P4jZZa7qja+uLZ8fppgofSsDTBGnUrAnNYrs1
XiFG7+jlohFkovWQOd81uFzynSPuhPXqBdpQ5vMLnzYRsRueD1ez1SktCbtJYb2a
6ylJzuJioIvNOwLsqkMs5bEm1V5C5XlcKXkpv4BDVOvcZW4YcDFCJbK5uOnEJdUI
dGqh7h6SOX8KwCf9z2RIvKmB4jJsq41gIjYgyW8Y9HXcwCMBD3PcHd6Oxvnqu7Ms
V9lrJDIyDLTYIEBTk/F3rV441C2Tit4TE+fcqNKqyK/pJW7FaWQVYQ//kIVWE7Sq
p9DlakOH+46BUUQf2S1eieakB58CF01lgmLu/g3UxrvtQSr1E1kIAwJCd56fg6tp
GbN0uRxWDWTCkxQZQZiM6/pqyYg8bpnRN5o9IlzvBWOQTRe+2x6qTdAdDKtF01si
ptvUUgMUNPnXSCmzldBm5nA/1srDq/4h/5pxaOAtXQEByVaZjsPysDh4sYcxtfl1
oI2md9lv90zoQeeOstKBDQef2WXDz3fO7SILgRUJPA6cgzUXKLTyZdfoY6QpCLP7
KajjJcJL5rfFM7TMjzXs1bhXguCiTabkejLLd447pLyDfE/0NfrShYr+Iy4ipxRI
Dxy83rxDRZ0h/2uwh+ri8LKgltsBtaap7n3ID3Pt9h2N5HJnUEO1df1pSyd7Bx9O
JnwWPv2hhQ3DK1k9OuzJEhzpICAquXRVFFpckqPrVIyGfFYU14Bhr0yjInOPUMM2
1nM6VN13OiMMzYtHxWrQosmOvFPtOtXAnpPNDQCtIsS95v2Z96wSXT/fd+BUom6t
vGcBhX/638c7TH87f0akFRFYQy48XXZGakepq97jm+c7ZZJtVGak7Sfx6kytiyOv
yJUhR1kyHxsIWbygHcZV2Of4oEnUgJgRtR4QDgikrBdnGIioFLF4Ko5e1SHguHu5
aSsK2vVBhHLM8hCL6rhDaR60oF8CIaO74cdyHjQ6OSLVEZx8sAzZq89smdAF0KTT
cExpoajXgWL7moo6pyG3JcSk+/U9q5+UhrNd0CWqsTt+BrEfaoL/zbizRKC/xEyz
C6S0tee7lmpI6dMFRBFscT06XowKm3E3zoT//HQQc1g3m9IuuaoBIJFe1GbXyEyT
hrJ5DPnHYlIfO/2OmHsdWORxYB1KD+EETcqxW8O/Xi57vottlUkyc7rOq0zJ8MOz
HQFok6WzMM83W+oogwQQ0DMfqnU5t+SDP43sfMXzYcuhidgGM0JE1nn69ybVbC/A
zh6EBoC6Q54K0fB0Dz5HJn1iphBfYh3k2HUdJsI+/MFGfeDWfpXlEoEdOP/sPKmI
BVmedRLcA7sqbz8K1LpXjo2uDV1UhQxzXmNnLoCjZ4UYpo9ysAC3uWkysca4mn8H
NXvgoYM7sOZSlZyKe9te8pyJh/B7vhIh+tYWhewNapJKmmfvCTWxPPSNG3VYXeSs
3BLJLxfH/I9mmOJnvkFkqCRkfcXyaKnYmTs+W9/CK4Pj+EPK9Xe2H+s9UWrrON0J
BUJ/QA9YmkLdzapssceoBcDAyuOmtHH9iLLhsfEOsgYKWdeKiTQYQMWwqcXXY2jU
6pakWuMxdiVXCAZLPRplHsTyMR3QslQXiXsxYYqbBLHbwjL97H1GTdT+D57zL/SE
nrZFIxFvBnxSgvjUm5Q55reWlIXKesmJNi+9e+2vizKcv+5OpoIU6JXIsTVY+xnx
1kSoqmbSF3WIU95trEsaC0HDMa88D9Pma/W2GvsyjD6V6bbE7OB+Pqlz91PmE+SI
uNkXgATWg7rY+lJQJ6j43fGcOr2v1/U1StFvqEDtAZs9Z5kQcgyQoOR57h1Icfl4
rizBh2gdCn1F3FypGFM0pF2kFQKGmzkufNNSjV0Y4bL9ON5GQwg7mH5BqfvHZN5q
RnsfcapNG+s8YkmkuNXIf5GyEei9wBeC5L7Z6zb3YllXWkC6Z9t0NiHOA3dpb1dt
eQmyhDZUrY+IdAKc44GEw14Vin0U/TcIklM54LrxhZf60+vsJwrTTxQ+QM+6JCD6
SdIESbBU67Vd0wsWhEKU34Bei2HzfpG5jyPnUugvLO8n/lxlT2lN8WbqKsYs0ewY
7WE9CX3rf0KrK6N9l0i5d1XVj/cc6lDGmRPCtmW4R8dxbm44qxSjyIofXzWWrUl/
HynHs190rTlmj2X5VQhiQDdHeWPlWS7wNEhpP0tK9dYiU4QE4FiyiY/0iyicbuOC
PatgyQ0v4tSHmyCh8deQ23EyjLkQZvX26PaPYxp65xjcUh8p8GvTCIhxy3togfL+
ZktatxWx0UeV9knQS0jGIz3uwVkrlD1X+aOVbR/2fdWMK71DfgkBCX6ptYkuZWsN
RNI4owwYszxqx9bz2T/YYu8K/XM6k+zZIUK6IPRAkr/K5TTPNu4PrJ/d76O7TiLC
rZnu0k3Lsu/4DFSA9FRxHKzVlWEIFY+JPntVbOqvpmVjSsQebN3F0Y79ugROFttn
CNveAL6SKFBYGJIUPzJ3C73A+g51/KkbUmqiASk2tNW1HN2bXLgIaRNkvzQtMmbj
1amqMjDD5nOPcjRQqWbkRCZUtceSvbQpE34kz6FNV5JYvvUL/22G+4NV0s3GX7Or
sVqU/vApfOkW+bEBJq9rdVLv+oPplB9RMwx/TeOZCFtbu8AnSzFHg5zEp5nWizUb
8VszbbYA4qfc8tD9kOPTKfePDFE5THPY6qFMwsHRptFAjooM5NikPOT6SEf74yZl
HvnSltwaDGWedY2c/etFV5wjQIbKkXgUPR2YJMGakm1LgmpNK9Ff9GHywRIz1lNd
2eqFfp777qRg9SjBvUtgsqYzkr/YTqI3bbvnjFyXpMXEgePFlfvq63+9RCdaiqGR
b6PxM/OtwdBsyRjWEaKW7JUn/FcQuhAzxSZpwjJkBP+KrPyMVhXHYOTPXxIDZIq9
f10IBpSv9pOQqcTzkwnUjJdufIA6B1LqTmJyiktA5PjWHxO155CD657YgSQsFmMP
ne2sp6CjRD59jYJQE3Om4FGCaVAaEfDME6+dByDNHHFHP4FTP74I5N08HW+0HQu2
Bf08rtfwmsGAYwFzbT6hbQTYlwQugFpWkhk4WEmN8aigdYZDTrB6/5EAwHopNQCh
6PgNOFTMFPpn6Rc+L3jXpFxh63jdByt/3LpLY/7FYXH+6ohNKQe2TiUKWtmHBZnQ
9DlSE/V86lqskof+MVtlX5KsYWPd21FhY8bv/rFAhH6tizBj4gJR5XsslLqipeYw
cpoZcDwIrPq6ZeaUE9Ui97MICd/foECnw1SQzmMU2XOhIAlxVjrXB6yy6AtIKhcD
8IsghytzXDoZXdgb6znsyIC0v1532eBq2E7zZOfjP0HhQ6X4NCzjiZLn+vkSQf3o
aOvdmvNlX7weVd+tMFFraOMcjyfeQhZ2zufUno22EPhFUC1Zxq0ehSP+zOo42Dca
BL9s/oFh0OdH7jOUV+5VhDS/h5vARDD5Awbv2Mu4gcd7w9vsz8AnlB5Z5Q2Pbpr1
upRPnO/QWjHmnadZ7NwcjQw7038s9FUi/8Buni2frs+4tzTbULlqFe7xfPiKToeo
oV6qQVOUqg/oMV11nwgJwBfWOK8jG/9efZBbCVjZJo5Ulh234tdWVczEbyX9Rjoe
JyRieE1N2dTEeO1xabcEYMtBKYJyKk+ettj+NATvnLG6JSrVRkhPvuLkyW46c9Dr
QgsHLloexUQii1yZNvLBwMN6wS12qXYFcYyGd9wa0dJiChr9m/FhKYbVeTpFSVP2
syYjuC+0HZs8l+pTTzxPC0V1N9DLQNXre/JJGS4lnfAzTVh/yo7Mlco9vVSxl9N9
Q+abfEn6SLLjqXjgpMDJykZkwpeAxiE7nwHOhvaGjB4DADQ8uRJmRdCHefT5Ps2/
/VDekIntM7CYDj96Ut/SHTUf1frhdtwXzJmSxk1Jp7Ip2K5BqgkWqC6wnj3WXyIQ
8H0AxPfI+a7yUNk1W20WSBzX866BVxMM7qNxqkauuMjrdhbO/p5ASW3kq5wWy8Ji
LRSml3eQ1QIDUl4Rdws+PbLahIJ+f4yWKHt33fJOIQ+d5M5cw+CYj5Y3kLY5E0aK
GvTW0nonVQ9n3Ss1EMBPmZxbj/PxWpsChjmBhhyPhH8b+FpxpSUlszPv5I9hBQIT
e+aV8ITrmGjR3cwLuuMl4ouC2lR+kF+lhdWDpqTnD0OAl+aZB4PrEnU6QxFbLQGU
rzcm/U2W3W2qZiheI16hFRJ18ACWURI8PjpoioLpMHENlSScd9NR6J5QDSj0seNJ
RASwPa83Ap3YvpIdl99yif9/9sU5ypN1Se2tJl022mKejapuOrTpB8qY7s8rhBIn
TUwR1VoutSPq0wbskwDAD44iiloaME7mF6AeTAFSwJJ3tSSsFBNU8OEITJVX1+h2
fyiyeZR10S+u4uemi9m45+1yjS0QBkObwFUifmxDbESDLndU88GM12VIUR0oK01D
YrrZOM0/vG/vV7VQQI1Q+YVb38/YkpxjCPk7yFvA00j0KmKYSS+WpaM5f8Qz47+d
1J1HsEbrVj/PBY8XlczPYI16PhTDIuTrLE74pwWQppgpqdg8PcGuNIJI7qMXmQl1
6VcwdQw4r0ovu8VgbtbeXCJPlUVpDLSh0rVfDbaNuzbs2OT3McsVZwjVon0BIiDE
4swJrMN5pAsEO7hoq6OhmkBcfSy06oTrvldp0ZmQReGHPCZ5KsJVqxc849DKzHq5
imeeBURYZaSCAbBZhjqKsa1fsG++VPhgKYhUbr1rbPoaWOmcSvojGhIaTIUL7+XH
nec6hiDE0brXjABpaeQyjweN0s8dPhMzMW4fXrTY55sg+KO8wsrNe0j2ErVdcg2T
ie/t2dl/A6LsOPUmo+WHbjtAZ85f+upPd9tFy46kMmbRuw+sybF9ZwR5eaAWrV1u
2Gpge5ZOTR2z0jxxdDsO+tIzlwzMxoH7HyNoZcXV073rNCynbtFnFahFlCsEgVAk
kn8dfLPIIqAWbcRo7n82rdFmbVL4bo4dNYPpt/PrSYVUyo+SuKjaBPlGdlG7V443
azgMnyC+5ZQoIqBaQI0etndjfaP5V+BHEowsd9c84uS6jkvq2XYcqlAza7H3SlRB
mbvIpFr5jCgu+GEsxPb1kWgCu7WFHHCfeUDQ8fkfcmtaNf47dTtVpO7Dg86S47f9
ZjsQoN0F5hffCUk1tZeeXAIKi/lagbBlTkWdCwHewLFg2/jJRU6LxLJQV+XYWlol
Q3+lnmP7QTrIrjLNSUhVBwKpX5d0aGaPtHJMdidepgOQN4E51TuSjhyGnK2iiAr1
N3tA8gMnHIQcBVX347fJyBN/jFhVQMlFeFe/N+5eW6LgBWO/ttGldZd6OQYLN2D8
Gb0SZOoF8u0tnDsOfR7BM0TeXc+7+F6XRzFFn6kRQIKs0xPfviXdRpBYoyFvfgPS
7pXiSYrH/KC7PfrFluOou4+2xD+OCAKrbeVcPli3v/E44j1W2vdKfzl+PZtMo3Xh
FRYXXSvwIjc1nR0aN9PEfVdWYpVIorIjHCf93yPiNNFJkB1B/Y4DBEHdD19Frcs5
U2pMQGiR5ta091unWEkJISh8MJPb1RRTQQmpjiuxVxnGI/cU6xgWM40FxZlYY/kU
algB0OHmjsUbef/kj3LQ9auZtTGNRe8xT9bXAy4PL3q46/8uRenWiEEZvVkaVhjd
M3+3cYv7as3pGKyBdrFfQkRnL4w9SDZivDdyl7ZJxCGJp7n1P51/kPf6M3rxOq8N
LJpMZezLg8xLP36Wqaiq6U1whenOKCXxXTVrFwEyG/gXXr0bc8KNDWU3dbQBaE7h
YGhQvSSw2+u1dNZ23N17ptBX8/kpshDO9SioCkVt9pJUKHgVWWHztA0qoXLqsNTz
hT+BY8+QqarDAPKH3r8PoTOkuxQt4SOJmvBqCVQz5Hk+D8DoBloQbr/wbSW6xeDQ
bkGHAa4+LiotAyDjU1PshxaLScRoaw8FQe5J1vD/EXoLgg1Xv0//USpbByowCuPt
yuAOLEx8aJFVuU0P+Hm+2cR3zaeiB0ejUIyxsyUSmd2XQtxUZSTNdrVMW0D1RSqO
beSIWS3jyi3AofcWUfHuL4mTKL0tBIqL91n9uaqyNZaDDyi+Vnf1J00XfLbk4pVj
MnMfpzLkst3ENMQIrF0p8EWxjiLSUkN/kQW6Og69qYnJKP0lqlOUQRf/ugYgZCLc
wIgk7ihs1d0ByNNGYj7b81oVAi5BK4D3gln+ZHOOb0cZz6ufIIRSSGD4MDfUUR9q
JvS8dXn9cdv5dl5himPYbdjfDAAjMm7ZmOuceKd0A+uqspXzy8u3iUmr9k4wNulA
C9q9y45RJbfhWYo/eSDPeC5vGQu/+WqHMApgxMUJz1+mEDBDQCjqGLbv45DVcQEm
sjtFPFRkcJS/5eX2D7pM4YiM0uTKvS7N3MERJKUYoV5p4d7V+WRIk7RNhzGGpEcO
66pycdNSaj33coILTZXfQl5CNWUg3rRqxI4zFOXlQkODYD0K1OMJZSBvDVXl3RXR
EIA9DxMIQbTiRkn3c0C7Q0zHzczoa3aLP1NoPC0YZFq6K877gcVl7/OC6ovvjt60
mOO5/l+wjdmnVm9cpZrNIyK48Xg3KM5ritHLYrTCteMLZGWO49y6MOzFDMWMldQS
VOxhAlxlvmacVKWX2yowZzLOLV9eAZ3tFugwmkwFCvkntdjcpDFkRw8slifdhuK0
sPa9f39ufC3NC7lIM/O6N6CR7g0tlATOK3fuO8tooXps8OREOQ0EnjuoY/03kWcX
Rf6RqNJi6ojN7E+09xETZtCP64jqtSMtPWvAl3s3uUgu1p1iU/bAl+vU95AMNeUA
jBgN0yfF3bN1z6lAikou//MP7Ewpv0voO3oSUCiLa+fgNxWDtqIcAYvsbWfEZQ4V
L/HFKSfFbiWvGT9y13gPJPcJVKMn5Zh35qkQL0WmstDZR5xfdWVqyZe75V+t3tS5
unzINlJJrhmewEffGF/HncC/itHt92sD9BzEAkDLgH2HIStK06A4z4EIcvpDJ+4o
Eq2NyVmBays/jkWAIk3YugkGUTsCpbMnmdFjLDcko2dUkrfOJkpiIgQ5CT7GiCaA
276Y4BGKL6dqV7n93gZBq/yZKf+p6JbTibkuHGL5QcL8lFi/TYGsTO2EryIpYNE8
NHvEYc7hmr3Mc1VRrRubC+/bGvAN4V+PSjpSNowDX0JF5lImMK0chrSnOItfO6Rz
yq/TDMiayonnOAIWBoYMUAPRWgsBHeb5XiYeKg0p5kvLa/AcUN5SsPA3LnNaoXRp
Z1HwBiB++2o4eTYp2ST/CzeTGgRMlp6bh9OAaXvfObccoJYDfnueNsA8nlsezG72
0ATMi5S6adxm4GOT+NctU3IvYEK2ADza8HqulYfedW2IPsb6AfqY22yp6QRia2XM
WVncQ1kpz4ee+knJX+TB70Hc8yOxvAy1iysVmsHGba/EpKjcunD5RVYbqGiAOUE/
aWZFblbXq8ke+ctNw6AdkPRDiNIH2KWtEIB1/qitQb71lniMB8rMKxynkdCPLime
pWuc++aEfZj1KwoJafi7hR00Xbg1vmywppSZTGFBGZAIsyMhZUCXBsMJUj/6h3F9
JkQwnM4/1AZWuxKai32sYO2+M1DFPISA7kVhzd36qDQDaU8ePbel0MxU1hNN5WbH
L0cS4D3VKFYYFSbjTrNG8laWLLZNpmsEWzE6jsN/dhkaID0kxZgMeiw09a8Z1foD
XTMwCgWEHtrKez8GBaBDbPOL2B9ZBfHV8+M57wyoutyuq4OKfEtH8puf6tadNr16
KcFD2uk0X1WbgPmrM0fGqt1J/ga690J8GdC6MFb9p3yLZl2l/wgINECK0L2L2Ixf
uwQikoQCD+RUT+RnxBnyjc9dn1LqibfIzApWKWhOp5x6LGzPuJ9V7qGyiV/JXgR4
PEQI42Um2nt1evZwPJQ76dd6/2Jmyp7+vrTZ8ZRJUcFsXQXoPCbxbe2mhZ97kYaA
4qWb3h/jMoQRsa7InthcsiapFijab17Z0ry0cpH1mVAvgLpIHxVzif9ur8+YBK8W
D0XRff32Vkx1v3E8exUNYnLWNE1rwWgIb1v2NMByTnDv3R7AkdaboYUhm+iNFFjl
MtXJlDmJUSIUV7AsnNdvkwCbckSunLEJR9VnoiBBN34suHB5Pij2H2xY9rPFE8wh
v+ROlw3jgCuvFCkcICQ+WAOplEelPs2+HscgD/gDML78qXuXhSem6ElLa/IYX0HD
TFOCxi1C3ydJnWs6NcYpTcD/PtDIq3wwH1tSGSEFPG8B+5hmhZBSEazS1tEwyhh3
aMtt9HlBrR3KAQIMv6Av6NfxIc/9JbgYJso3LMNsQXhpetmwdtVodWP4ALhRAYBc
4g27y8dXZP6pGs6fmATcHUTVskJLsiV4BWqEzJNfmqwrDAcTMZxapOhlHVs6UP+y
wbZJODQGjS5jOa7PbVz5/vY41XesivUirzY9F3hcZ5SejNiBGzvujJqrCZQycNty
yKu8/JBQWT3NmZQS7goH3FdS/sZAucMqSXB7U3SsuUlxLWGVLqhJ2tiV66kqYE4v
6bA4uD91HXkJNCwOdLa6kRZh5svFOPUqo1UfiUmmdDab6hL9wvjAYuQ5g2NPUzGS
N1O3H9aGs84iIFp/G1Vc0h5PsuYlOz5ybNF1K4KzfZBfweVL9601k5c+IrURG/6S
UWU/0qd3Z00+ruan1ZjBb4jRS4reVtWG5QJhC7J975GAWUJPhibGWcK+pR0oF424
SSKma1Eqw8X14QMPIGJNRIjTYjpLXE9z+K7lL6DPs71FAwPlih7/t5xzNA4FSKbZ
Y2lI68gbjDhO13vSC1UpocIucujuFBVpWa7Y8AvfYcOnEZ/qtuM08XwRTOuEYA09
vSLlh3k89hiKEfIdUB24NxiUZrjhyuEpIeAVD65PvAwUq4PpHkI4LNayGiwhzbYV
tVd4QBl2teOa0OlM02IzlmQhzgjuVIiKJ2Ki+aUTn/D6xRhJkheknZYj6vEHktqG
RMXYMcW3QiMkBFW7Ijw0vvXfTwgoH6jpS3o42fCAK8PJ4Ty2MhVTlEXET6lY1iV5
L0VeKAg6DIXu0gj5ufc57LylsUyUGrIDB9BCBaBYyCEwVuK/DPANKxuIVIuP1gjg
6GKO8Nla5DKWmbtV+g7xmA9x9LhlMHoU1exIjy3SVhqeWKTgdWgDiJ3gvQ41i2KW
Zk5wXQWwSlSJogrYCrdUqnqQ9/kFj28pSN1c9NcfC7B1wl+gN1K31xqzos6Py66D
s/KfNObmGGP9SWhwuBztVb23fNsQZfvcKMt3Dz3+OiBHLCjA61nQ1qgmlbYQ6Lxm
cJvkKsHGr4QbWEG3zMl9aqRhjOdZVt+ZOcDXlROrhsaAdavrBd5O0pCwZO+O8ZcF
wgpUQ+fkKY6F77nWE88R0b9SJSKuOCSPI7LlR48e1cgOjPEFJeR24CgZPzJHOWET
pVpEiy4Kl29NuT5dyyHenMDsPol0YIvRcyK7rDY8rCSKhjCsB52Q3zqXkiU5MBzc
GsOHnB3D9d9t448VD15gLdnx5t0xOf0epaGHTK0mgI88MJd31WO4VqS1QsOSd5Y0
7e6SW4ouIxJxFeFxeKg1di7HDBZeZps9gZ85BqxwRPMyFSxaQ44MgII7D+jKIJZS
fYGaE3WJx2tRyCYBeOeuceNd5rBVpsUuKTqGV411zeHvx4S1xrBLm3CChgf2kzRj
/WTRwqD06XUWSEakvzhlKlSKyZGTRMYMrEeau+ckzm+Xxz388Rx5LB+KbwByMlD3
AMkt0PcsoYSj5b8yx6l3mInIgiRmC1Ob4rJcmxWADHA4eDahhPZGbKeyyrOkcFgL
qXCS0ofOSHiL1zxLJm5KOlvNm2wLktGFJF0ehjyBayOQXrnWRvsAkxPPECexjWLh
7QYlNvN//qaFdF+3bdM674LH6zxgiCgL9TF6v8PPLo0wrhcpX8qWaxRVweESgE5v
tx4VoL85veyLWbxBJS++4agoTTWvt8wOsvCV2+7M+g0OEaeRL6pv5IBwdsJo3dTS
3w1PJ1/renXDMhHqwY3gX6nfqAbde4Xw7IiylVwCnGQUaXJjl2uHAw871lkN/1Ea
sSKve94jDk9VfBB3SK4xT5KBMHSALtY+0GFnqIvGtHg4LtTbSgGuVth09DrSoDpM
Ezama6ypyYqFM46gKcuO9e8xPkQGUV4Hx9E4QmsauVvX1moPKddtj9KWj0mp1xZ8
Ip7GA8VY7Ph5LluEkNBO7CK/Cz5WWm9eI2czgbCE/c63TTFQ+wkGfkiPampxOgAI
8753aVn0kBP0khkaptavNoXHVmgEVY4YyY8HfaLaPW34GALSoxr0/jjRb1Y6jHxU
zicRkTzi7MJCxJ48QqGhQr0KjlJbD80XEM7XncNFPb96v4I382eTiPQPthCIaXN2
mGh+IxiS5Hy/BNSLPA4G6a9PmRKyl8Okn75+LZKjuwSk6+wu6lbIbXkNn2klHnWf
QI12mEO0Tg/eXI77xlcr+BJLJlV58PSLrKNyZ+iQKA8k9qwAMlT03G79rCYYnRnR
rHZ16/sQibE0EO4mjHdZ7efqPn2Of1O3/nw7joMtfDb1LTTzpTNDRCSTgyy4Pp7H
87PKVh168bmNs61If5VEJbLphwsKIHPEo4phrXWo78tB86OQVcwpd+tjDqRaWkyY
daub4heD2UWQ6cN/urw0I4Kouu5jmPBNkW57mb3qiFpS2HjsTw7s/LiEfjKd4KBG
T0TmBeKbMTFECm7+NwGFIV8fMUxk4e/8uuARZsMeTXEeBa1w4/yPVu2EPkTX+Y4M
0rJljB4IFAc+imiCNfIXNBEkuFDRYDBSUWno6BxLo/821iDth08FHEEdtcp1Boji
R066F5t8CataH4A0JpIvQ7SEv0sqsFCo3i7YNBxUEAMD0syXFaVKk4A2jF70gyqb
zQq+zsjY/KU3MakGA1LoPA8i5XOVNYaeFMlPC/rCWNk6uaVRSh7bvjdDIkJxEYHk
voDwW7Qmv57VuB5d3vSL1YC8iQSfWqn++eSW2QuaEyD1moyxAzQNRraLa7MZKeml
aG9gZIOuD2RF1uAQqLbWDAtSj9XASszn9T3L0ucz2XdwnfI3RZURnoEHAS9YKvXW
WklX4ESatLMPUaAmZhXgaUZFaqlxS/jAEquzvASnglb2n5Wq499l9RZmkFTkT0ZZ
36udfhvWuoBc6/xtvtUCD3rtkXpQFse/BMEr1JCMj40g1WTI2kbwJkyB0+bhEnao
MARyWbSP2xOQ0CPNH+LA1zjQ4L9KPeEZHS8sMDXRoczRgT5Yg4ZEaqFkYhVkx9xa
FDEctdLxHWczo4U+Hsy4R6kPfxOgpv5MNorlHrLSLjJaHenNy3aCzA6hHtdqxfP3
KucVq/Ii1oQ6bEBaFHP1FpU8IFjLmUo7eSuPybJQ9le5esj51f1thSwebwcUca1I
BQGRioGBzHVz8eO3HK474Im9mfiRD5EClSOPnCxQ8MA63uR9ykwyNbzWV03lP9Lw
rtkd640RpBFOFy7e/JoXdhM6JMuvyssGEe4x+vLFsp4JTi7+z8wBmF3E/wKj+cTy
oYtlQpxnZKmTJfo2L1wCa9mLwTcPTSkSqMyP2SvpOHQBpAkM32Ouo4xKwZJ9zQvL
dSb6kaKG9LF8NJy+yAlz5E4tL11zM1Kjsr0fshCtwZpUDoK+fEbp048e+Vz+MsdT
OpShZF7wo5NM6DHdkmuF1OyN7fU2KGerUBzdVniZEzXiIbB/NtAVgQtthGIZAzC7
lu2vR6+lrTgqhJLj/UlhFbS/RbMuwAXmzeTnd9IBoPt0/Y2An+OmVLAOPqEcAC/P
O44RIrtsaADM8V9AslMi5SdLXPan0AzCFm+R7xDaSDjwKD3hNt1OXh3NF7mmCdZP
ABKEINhBxzY5SPfpNKE3Rl3jfqsdCSe8f8mS/zZq0CbYBWFJmqvWdM1D5r4A2Zmx
exkNUQkWlvSK7sORtHa2RfvjfEuJ8OFbdAZBMFjgq1MQuEk823CvMTJXKXPi8uGO
0cGfj6Q/KkeXzx16qaiHebjqY2jfDEutr4/aBS+FbothhRb5uXBMsqvnK/ga+CfB
F/IIWvG0CGNQSgslR+Qnt928q6A/5WN+b3rwaipW9gGyRAJlX7APhVNgq8MpBbQq
cB+hrT4oN6Rj/eFqA7o0JY2zI+lzrgedZ8HxNoG3m+stZyNc5nCKoPWZ4hnaR33z
mfMcYSISth2kOuk6OLNbzJxiORAnj1Vxq7Pqh2GAPcC1iAEE9tMyA+WnhKw2Ibts
GhiGKNnuijUoMFOPdvnU0bJQYRLQTfdTSfaYtLQW1hYldwGRyfdIcGkALXz4Or2D
mhGC/LYfvl1MAMu3St36LnszjVXDBIcEyUixAtawnyNdUi8wGq5XxQLTDbGyq4J1
zmgqy7hI9LPURJv8hnDU5mn3IwnEaaf5H+Qymrf+dAvuuy6RBeTYiEHiXxeZANiP
AScHZ/ACP2i/uBj8YuThgYJNI214uIvJIY8XWGNnRtQ/RZW+OLZtf3T2vWCF7mwQ
OVI3/gVpHes7IeI2He8211zGeKZpYhnvhEW+ZYg2C0wxKwrp60xeTiNX8DJuMKl+
fR6Lbf3j0GfE8sllifSUJhauUafeSp7YEQpfazbwGayaC9CJ1lNmP1fo7ZEUuTSZ
twdnPu9c4J6VqoBhHBx5qkKFbhxzukebSlFYL8qtiFnMRYhWhQdXS7c3/xCIAPbG
IhiuZYjUjXf88uEi5Ek447Uq3R7kSt/8CVDEr67FAFkqD5j/Knu4q99fNTuoAckL
t1wYzwLz2823+rJgNs0TSkl8RnFFw1vlQcMzc4yBoJpusbOro3U7a4qQHZtKwKRo
POAJ5W5Uz0sy6JKNGMaaVFziEUOesHVUPZK2X9/1BiXvSG79AEVK98Eg13hc9A6k
7EdLwtTCiQOuJHh62wsxJVMjvQm5H0JYlALmAA8eCZfxGaQXXVw8HyAPFpjCKAwu
hesUmPyoIT5HSjNx1mseWRLUHMFkfigi9rDQoIZdeJfJdl5CevWCRYdYMGWCuZLv
+Iqu10nXPdcBzkekIIKod1x/o+t1OrBDz73BpqE8NmVFqmrWO10zPK9JSPkFaF8A
3TPdnHCqFvryb2+tQ4ip7dO6zWC56bIuDKaoRYT5e4ME48N1gSV49M8nG1FYpuHA
u9O6hOtIKgQxaK0+tn8vO2Htv5t1bNzc65KLBq2Oifl4TKivTRuGU4mj49IWqcWj
Mho3tT+1w4/WA1rdwOhgzJlVjHB7TwpqhuHLP+FRDASz+TRAGSl8J9Rg7PD2TaTd
A1zFS6YIXhgTu+4QT0t/3pM/4DDDuqtad2an74aHeMlmJ6tOIHJr/k0lISH9ToTY
vzAO/nsflJ+nATSmhwBj4drjT51AHMFFHrudLDBLE+Fa+f7kY60WUOobnvb0h+/e
9zQIihxhv92erQhCiDJ/CT6vIiiQV9Eepv/y5QTP2WWeBKuE+aN0Qs7B6tFbx3ZQ
ArU8TnYYeYIIUeIFeTTsSdmiUFqVO6SQ4u7whARPYJaaXm7dVQqxFKmPlazorOdZ
LlJ5UuBn/QdeN6dHVTW1D/kSDK5R4Z7q4ib02qnzqGm4qhGESWvY9klNthyg+pFa
YlxvzfSnh7bZalamUHHJ3RE/80I+SNnpRA3Dt620ACwbIpCSOSaCMVRdlGxpSmdq
rF4JGjtfPsFHm7tUrLXCcqoUOKZw9qtKpkAJEreQDFay5H5tlkvnu7vqRbKrLlco
jm/Q8DrwcBXWCu9ATlOOP818iAlnuihzc+IgJUkl4z41UAiVl96Hx8fxUq3Y7VTa
m7W/mCjmKpiqxi3NjgYUDFGd79TiYn/Ixr5rgPhHd7yi05ToKF3nc0V20hlDrsHd
4sf2nfiKYtdQDRh7+p/tfL8WWGe6bJKVxPsR6UtKaqb9JoMpj3VG7u/pjYsAsRJV
iSrBw178MDeBf/r4IyzC0HJ/a0wXKAoEYQeqpu/9lHeO/1lwpYa9L4wsE8Rydbri
i1fMn3lJRniiHPytcjcsD0fP88WIG3/l1A8F+oZ/+nM5ArmCXu0ZYxTdVz+zQ3us
L0zR1fdirCnXC/77Q2Ha8d2s5UK8iecHK/ogtYp9KhV4K9IoCsVIjR6r3nNZULM/
iK9ovc36i0fSkppUjQ5mR6CpD4iqM2pZHJ3/eGubTJC7Yrjf9zucPCG1N+rxBKcW
eWmrwC4Bc64dl43JWnUqFUT1tIHlsGzBAzY5Pl8MId79+0tZir7ivxAqu4UeuNwK
nff0B73Z6X+xolrsDHZ+2adJLvVsX4npq9Tafj9u96bMflAX2EUdGfdZ+qqRT79N
gzhzT3O3EVGaq1ZRRzf7lfqUMb6P94LEgcHMl8Nu0fopyorVm/5FWPnIE5dG45rz
idDZD1KNdOspDSnC/12bdl/g0z6oz4bHnzJExuV//py0B5SuDcV1sk1nFPu8IgPC
Ow99XViCs0pFlS8HUBIX8/AwmtmMSGkV7w/pEwlNAlgjtZedSlOu9NG84mBa3Hao
Ute4CLUYz9v/abO7FvOybyEpqNSmkfNGg1Ayyldm1FDEJy/lVj31998ov8VjhTqW
SFscJvpf0PN3CSIxWfgfrVIS1Z9y6vEJndGAj1IXGogfaqUhT+1mrf37fybgZIue
IsuWX23lDWZJ+or4SMBUUrjASSofhxsE01ho3bCNs400PrtTvTeMB89n1Kayhbjf
eEwR83oGVmpFt7XoX+vg582juGOIAPmm+7xR6CSv4r/ryvNmeEwddkr2LQbElzKj
jt8szjy5TMiWqO88z1uZY3IY4o4t9K8TQGWCD5fv+kI0njWzHek8KXmxyT6xiouc
157aLggoaUkoPbYzMnsVOtCjZ8MVXKRw5W5zHj5IJGukyFJpGvCz2WTOtRM4rqn/
JsmZBNvsWVITkR4PUnoksTBIFHxMsrh61cCbmtWAXBWt85nw50v2GFQtbOL1lCBE
HxHdmKOl+Ne3m9SKDvC+8Vi2vMUIuhUhSzjfvBgVyCIJhy3dlfbPYGCSsp6UwBMk
vdXDtuowSy42bu4BRoitVm9gTHqh/rm5W2OO1rXTNeY9GDnQUqR19WPt/7Wx5gyB
zB8xoqctsblE2dHlxiV89Ju9h8iUIPpetSwrwWc9UHhUVJPSDJh606bEwr+k0qkf
7sg7bVml2kbobhhfrfr8NToGxGztJNdkWgFE9nlJbZh4nAqbTxiO5H/yZDQ77ufY
5iQchk4MYkyXqBjDggnre4yityHUsNgAn83GhPlOzdCLCkYY4pVMKcm1Q8OAmp9C
KP/8DwXa+V/RJOwenauanpyJj01wPG4vp899CbXao+JzrMambeGmxX1XLiWLCB5e
S2y7sDkNHuGn3RBEXL2pNgZkdirFwKeafGsZaFhIUW5FWllqHir2c8DpWLca/J1p
3PY/Spa69w/1PBPkPVIpGTJxHec0NPy6mptz4YlVe8bblICLoQCh8esb8lvT3nZ5
FCppHeYQrYCuUCH3VWd+PT0k8XBbvFoxo7J9qr7qnRr47F5py1AKVJ0M9Goe+S24
eVRwmM9cs7s7kbSrvyn4p3B9IJoihiUXwY14GtBKAfWO4MJtaSMa/+j6JuYX0b0t
CCWzdmd5JujCPtprJtzRY6/q3kYY6PAxZG0pAGoJZhWsqXgIqCVVQX7mzKzJL1Ed
fkgnptSvD78TaZYbMDOKlbnOVefma+I4F7y0pIiwwj7shxTTob4eoARFwywmkI5u
5JMO8NZqoeEV/dpy9hnxDCeA1J9rMLnTAczhh3oPE0Qi7FQdyOe6nm3hYbbnjvs0
/wViY3eQgK4i3X5kCaFpaclDiWAn56+uRAEkMXGCG7LHT0q74Vm/sZjY+Qj080Im
A+fbDNi0QpQiJeKQFU+FLjnbbep++xQ3xmR6CXPN7Us/cNYy5p6lSTiCZPHLThX/
be7f8EuHcA5+HE6Pn4HY9RQK7fj88bBbV2+3GDQanJs4rbfyFKQUEKCDOP4kW0z+
lZ8szoVPuPhqbPOm+lSwMcYW4ZK7/UaJbMsLXfYwFUSjH78wgqiTc8HNFQV+K2Dg
CUzGFgHyS86zTrbtVTwiuQtQ98wmMLqKXmEXRwZF7EAJ/SNYpNNfRVNxK03Oeq/6
YiLC+FElxol4yl8dNkJ34PmehJAqtqQyhgvIdA4yEK7GPhiWLdqPxIEUNCE2KTFb
qooiWXWW8FMP2w9HDdu5nWWNdGq4aBuBw+zrj9qYAjgoDVpR6mOPFDdelpHs/rUy
EcAX39kiV3+XoTDplaLEN6EqiEZv+PX0oyJIK1EEU6s+CcN1oiqe2vUTXBbNAZMs
qkMFiV836UwnbNPv02urp5chmrhSo6Ees2GAXIbxJvL2NpQpJD0jkQ18rHtuxWWi
0VSbKUxygT2+CAhTHVNBUq2lBGmXR1/xJypjnHYYtGBj7ec+cDi4MipzBh/mNl3w
vPvzN+YS58WfOARFiQ6fKIPWRcWqOewb7U90MIoAsSb7xOGhNT4AoRZpPdjL0wRg
Tiygb03aA4uJOr5YDidGqiyaTjGB6NDDG52ZEd4l3XYwQAUS1CTDs2XJWHVVl4io
gg0a/cYZWweUwaRTWReCb5SJnjAj57XXt+7XhO0fykRBkz4IWJ6ymaY31Asg/MoN
G5k8xe49K0n+PgeI0ZwZsj2OOT1400zDtgw8rghPTN51uqGBDeUdzUsb1BMqvLV6
dg7cTaYiw+K0SjN65iarQOmtHmlf+Zu3arIWNf/+L92UEjIIoYo7Dsjh6m0G2AFz
2Bq1IInlyBbOE1gML78f2Y1Q0uxb+lprjbAFZ3CcnO6eZQyiuHwSPqq3v4pq2wbU
HyUCXH8DOcdlLbukXVeEmGeoDN3kXr0YjoDNBwjfYMui8ztGed7hdRLWGyMnf2VZ
J+gMnZEEpMjuAf1ObMYehEurB224QyE6h9LOYjqF6a2dQUbCra64bu8e46TOwJnF
XzU3h0uk0feedk71rpqFPXdV8/pgnnXYXyWpEK0qG2vHTRGYXTSb3wLKjLORXZVC
9woUwfPsoSlL0h9BAcEHaN39CZw8Tt3eoSgipYjUDMbpL9WVOHA41QCBQx5KBT9V
QtjcdRf8KVSPNO3b1TNPndUepznR+2EyrZZfOhEADyLosKbmljhot3AmsYTNIfee
jSUFjxVXrtDEqj1IEN7WDizFlywrpbGVgmWvdAG3d4W3suVXowwPCVIvGUdrTFUN
xGqk8I9fHSRns+YTJm9WT4tT191ywuvv2IwW6Cl6TU0K70JjFjPVRHsp0scd2KWh
DKzyOr4Au5zD2nncyq3j/J2FsBGJdRKWyp9sHPc9D3sw5K9RU076xoroHqvZoz/p
TeEKLo3JoAXJ/S3KX3vHXqwG3jlJWldpRWhtl+H73r4HRIPK3wgeW09UepMoBKW9
Nv+1WGzfT7PNnFYiA2SHcrxKHnhwGb0FSaMpUMID8KJ9mrxYU7eW/hdcxm1fpZF5
Ek2erWDQw5mPSPX3InQtZArncbzN1VqnuZ0vfxGDwL0JzbpODYuYWCZmYwm4avEX
hsxbIyUDH6jYNJyXVUOyE13lEI6A4B9d89mmN18BESXvOzYm8ddKqCeqPYfpEhtf
CgXn8yz1SmmPZNh3YlBjihGRDG4QXSGhlhEJ4XgQ4IwkJEeSyEo9QeC8nsNYPiro
bRS6XVXdoFpQyObtaXI22W74REctDM6v6AZHJ/CgOqBG4oXKyLP9hE/1goqz9u73
zv0XXtJS1NYwIQNKxx0pyuW3OiAX7CxabpvT5M0jFMiWxsj4wYcZHcto6UvTtEqu
E6onQtbrqFRRp4bG6K3hbkvrtCi3pbjSq4lxQ96lOlyzr6khrJQ3sKDGfs4M7c+Z
Qnch3yRJQ++7LQT4RsETaBydiY65aLXzxByTls3F43lFkxXvZLnukUVKbzaZC6SL
zgmlYtwT4Ko85OstwMtffHnLXt42BjlxmJjVbQYOGhwiYDBZYTnV2YPs+L3oxYxS
gudTEdLZXtc3vzdFoUg99YcKMuzKEQlY023jvgslSOHOoKmvwpRtAtd7RHAcfHxc
2MC1kRq0B6BrQAPVxs11a/fODaI855EmPvaTyXEPORd2YSkNB7/TZv3zovSUzZ0z
QHwatQ2FA73nQXnLYOe4uFb8W3euuhLx2A2aQoNw9+Z18IV+JKl4WnqnVaV1Yhyd
vL7U/Umts3nOj09MXWVq+YI0zVXY2lNe2GXQhqbfMwkovZC7RTnkow2flo3yOnFm
LSC9awh/Bz3OyBCSl6BaaEDVftBTcD4goSZb2bGRXBazIBibq615h6tCXEu/fHau
vtdxPKgQyJMnl/V+7srWPpYKNImZZJ0gx6pepGce89QKkJHFKJ2kSWHTBw/JgDet
sHHKwqNj4X2sTx0lTaLN54rvYdZC1IWcfFMYj/lS+5ItLdAEwz7pyUY/Mjtcs09D
i5g01hsfFp+PF7WhglaSZ7AEn/u6C8pY/HX2XtzUTHZWsRPy4ocb70C4zhZxKBhW
bJI7CS+RGfYg+f/aUMp8zxBq7W8B6YlsdmRrytvGc/HoknDOjqt72clS0Nni0C3t
rwC46zn+ooiNSAjjugvcjxQ61djR/QiaHKsd/ylPSwnxCLNsQD8/mWlpIP+X6ckC
4xCCviFPjsjG7N66dy61UQeSQCOfWR0q1YJp7Rn4/QLp1mdd56FZP01LxkVccc0E
77i81BQjpat6OV9GP+s5+FDiYnULT/aKB2WaJMyt0mABAYKbbNy7eNt/Jk7gzKNX
ccLoNzKlRAXuaU/gMBv+9Qtk1lWu5JlYHdbiGayvQqrQds3jMcX3I6dh6M6GYVRb
xaZT9sFO52tbMoOo/ps5RpjH9mMbUGBVyBsoRMx+/up3d/3Y6gpx5KjD01WgKX2K
rph45tEMtYIt0/B09UNrvy2tOgRBdQl81onjnlToGB3mVzQP/iPuxZKgsDz7jSG+
IpvS9Imw6WTmYf1U0oXqFZEVcKANzTA2TNUgFItcIPpHxPnrh9HWsHpe7ybMxFKD
NOr8x68GP0qd8BLKUViNoP/bQTahA+fTAIk7PxHxUuc/MukGFu34MmoYMnRsrfXl
37/X9YPm+q5QTIrepWUMFhkBIk1lZiUJwKa+e8Uu17E8mq6nD4aC6IiZdDbXeGVI
KFlDbIAWmuymOhNqwAK7B/g3ncikup24OoTSUB7bLHzvXzBA3cJzGCdvGdyerzzy
EY5RI2o/kkSyBZPiH5i3QBxtZBWKztGw45/FXqW3A2wHi9HFRn6JpsVsYL1z/vTG
3+uZKbAooR2QZ7cEm8rB3pENdCpgFzVwPIFfHtLas8vl1K+Y1drg5sXOpqz4v12x
iU4sMgj1EKDoyZ31JPFSG7rsnE0xhWwsNTK7nYYt6fqv7sjQQtj3A6009oDNXOSE
1u1n433mk83UfNaLd+k04CmG2lrCLmASplicf48AnyCAuMCfzzsIMcq7JSGAsQBj
Z9lBizK627LuWUv9wYhS8E7yCe+0lRgZ/N3SWTqYsvy4BvoIfDtc44LOlpMyiCQY
qvvPWIVPs0DNKbMxbkVtnU4v4k3HqAB6ZMjl40p/mw2mIy2wMQy89CcXo5HCv85V
mJQnPqlgcXIJ4a+NXFSYtTYscoUJY2Z9cuHkVBMACeATR5ywoZewEMXXXfdL7B47
inyH7TFS2ryr19BlMCs+1r4foGWn/VB1CKPXR6rKLkB9r0QNj3ek5LukGH5Y9gt/
LBVPDNwxuwqZvXNY3onXsieLOUeJMVo5PF5c2AX096aIWWh2/6zUCra5m8Id/PTo
5MsZUqcHFuTNz/F4p4E89n5uiHo34eB1Y7qsc5bDVy4kWhZIOnzoFLa/942p128Y
Tsl/KfO7vMJ/1eL3KlgJCzdFY/lg78WFgQWSShOIcsJSryLmYtegZJFxHfYvScB5
IEeu5ciUQekAVEYtbAhhf08kkhNhBlLdQRx2bWAmuhHN6Rd64z5c6Gl9j3oanWBX
oavD+WnTD8A7qPzzG279rEG13BaOqZMQaUvrXHkMnuL/+FtDSn4BU1VWltUgItNj
f62RDSj/xGL8WJ0ej2ZxYd9lP08uB7roubn6oYsVmlxniiEU8cqnyZn+1e7bqIXP
FEqAc8Avk4ru0akyUt3CCYNx82XZRsBFPk/Dor1y/CXaXJ5ZYjRawVvIzpitzx97
b5QP5s7aQQR1ZAhsbSESvKURTSMLEJKvu0mFoTJn32iAXslv2pvWvCOJH+7cvmf5
tat4zMPBHKT5UFfWBpkC6u9UWyH3FWFxUuHmmimuTxz5m2RvQ+RGd3cEQEujbJ3S
JukQdM93LzzWcObt/5RQYAcZeSF3i5od9ZgSEaa33uQ1OsfKxiLlne1SZ9/iG+4Z
4EYVrL6LVPO/nFYRtp9eTvepVMEIkGs6ndH+tCPEmW2cLhOOpxjMpInaVfebBip2
FE7stAxgq4UsU1b5wMdPymZUGVctFD7gKE7FKNkUYvXTgzNryi+9McG2ZiTH1xMh
Wbdc9ipsorPJa4QwOVQt8OnV6U3f24micoOjJxOEkwMtQBZdfsqplNJertJYXkQX
x00xKsHvskPB7sGsnxdrcM+Fz5Xe4HoJV31DnWWC5/R1sEFs+9Oy+kY1h+DdeW3O
XMDAlhWYcuGt2cge8ieGbQLniUfP70rBFsyauVa1YOUR59aoDSjfQxTtqY59IrHr
O+ww/iHH0N1dcKSNV3NtUym9IP8Jz1T/GteVWisi3OMw3hMy06fRVFbW591zk0yv
oZZzq+8+rjvtDXXeiOBI/CZK7FoXvDLMmrqy62oBJaurnE2orWKzVrwsV8+fJPIj
Jrx4Y73smItDvB//MPLJstFtqOg6ZfFpGa0mR+LmOOZyoV2YHpEbV4VD+GoacYVg
+OyWshoR/kd84PfcVutDiHDO0dLLwWS3C9+fc2xd2x02dc823r/CxIn8nO3sOdNq
lAsTbQdzayKCErucVlTcaoscyJecwu3bxIug2gcawq4ACQ/Fa+kXeHlgiVhWJDv8
Y0PyhnS+oQw0wBl+xzvEnlkH7L6EGlTwtlEH2hkpTqGJ0MyYsuOSdhs5Ap+VchiX
0IORBgDGREBGS3eBbLZ3LIyBtYRKGdAxemZSSaRQ/ka+RszBi1PmOeMVUi4tK79N
/fcHZZQPcrXsqlgUNRGNx/OaIRF0iQXWEVkKwXafnZuf3BFNHEmagBz6rfUkw3eS
XPQYDgVoYXY7gtPzwjOdZf478S7CIptIlxdsS5ZA2t0jiQFrGGdjEM95+tzRduho
M4bsrK/driUholD5SJvgg6X/9aOyEXVX2vVsM+J0QlOR82SVl9+tIvP9bnS1o5No
+jaAn33GTks+f1RuLLc3RHby0nkDdAcg4uhkhwIlrP0cPjf8+9RNQ2uq+Fy0XNN2
f8fvN7X9gFebQ7q89h0wh56q6Q1yykdDGhCJYAWDxqxfl9turfSyVFlZb7ZotCTU
7VqmpholqEwI/K2qbJiddZA3xAPa2R6p46dzsTAEhmIWfg+KcepJC6hZJ5k9wCWz
tRDL4kIUvO6QqpvL/lF0y8R6dN1p5/o+z2OVxRV3ouN2rVkStTykqfzb2GYGcRHT
eAKqYpVxsiUpM2khjLuNdjrpVm7VS+TVp8vMuaPfKBS8pnPnouHySZAv8O7FkHYp
JxbAsRc4krTk0EyyM+Lc8yhiMozMxVpQTfXoY1BnxAsApIE8RU71qo6QpHjTukh8
3WUL4akwhyP9HwOZkVA2MV8DAA0BOyNKNEN1EYGf2CxvrQfPbhZDpL9BJ5JesrNQ
TmXMvgQg29kSaxm5Y5atXlWhhpmtBuyRgBFEcH3rpqXs+H3rdd7sl6GZ7CeWUnIY
2A+MZl/asO1tUEL8T5hDyjr6JZmM6hk0mASl8vwJPUZVSk8X0Tg9+g75oqBo3Ie4
KVTGZj/v+yEexji4TwXVVgQEYgmGjKq9lqLju/A7Iiet0BYy5QA4RNyNjcMQS/gU
aUESUt4wpI3ijQZvG5hLHyq2graPl+NOMR6Y65RZMfVTfdw/YZTeTJRyNs4ZpLK3
pwzx5LjyUdYsdHts2dhqEo8fVTXiZyNLCfus062EQ9VYoZT4vU04JgdnPvef0Tti
nJI1bUqm6QvpXeBKli+FpUKEjvbMCJgm6QRTvezcPkK7D0+DYezHQozYSaD8N7E7
F/hXkL98fHrWKJbPQRcNejj/lRGiEyG5iVCPLGtvILEJZbLpxvS/56iNfZgl9BWe
JQb0xvU1SEOv4r80dj0n/dw1l2pvHSpFMDB9oSamhCnCR17yQFh/ShXGaDe/gELu
WMbTk0J+Ekg3uCndCHPJfEVKibIGxXaW2xmTIDLh41lImG59F6OEOZErkoXJEA8q
ZnXOH7wCfYLmV5jw6O/N3s19V6ZdEQoUNmwHDSgfEn2ext0ftD/XAIopgdse6Rom
0KLdyq5DD4xUrMRoxjzyuqQIBKLFLRVVdHrtXt/E9Owz5T1NZ7XBYujB0tp3eGqz
j//frhTA9o7v/P8nWhSpakpLTBnr9E2og9fNtnYY6Qku48otkO5o2GpKOC4ldUE9
T6Vt25HO5jE17bdhj5/kV3uTigVUqAmlC3StkoflD3+KhsiCWINw5A2AzNtRv+lu
vFDsiZg/j5MBTdWbeS+dqHteORJFEHfhgdmofOOXI0j5HW77IIwhO0pKcSCrAJq2
cnp9fPDaj1j9Di4mXKp7YXPJxtJGYQEusa50dcXjTKCUu+57q1wdJQOa/EKIB2/Y
Y4gMCd0MoKbgIZ1jctMRw/niq4V+11GxxuNjEXbzkAES1DwKC+R6AvRBhjalF4Hc
Hx3uzmpXBuSRLRmGzPKUeuLSd4qbPqTl1bNNl7vEsYldI11NLKjm7td/G7ouyFK3
gWHdHznsyWekaaKpMx8BB/sPECcbOt3/Y0Igx1mGez5TAb3Davph5bWjfecO8b6n
Un88AZRAs7UrHv5GnEYV3dzY3QMeyhzLZKxqQ07HrPDn3yE1xe7nA/BuulG1YHsU
EnrM0hbde2uLMJaqTI76nN73TRln2LxJBW76WMoiDThdr0sPKZOPVYiqV+gGQ0VL
LlxI5Q+sHwRlFqVJnyXftS3VBtAhoYSjszM1A2p17pZm7SiaY5qB3kg/1x0Phs3S
Ay3CwwuYCT1SRszNNun6Q4nhssPmruW9pwHh1N7EDgPqYLE3DoDq73/ebjHTL/6+
m47UaLIN/Ej0rpZ9klChJg+cTY0LK0eL6lqZbfSuVS2a+lcwI+cuNLK1h4xQaCha
1tO1RUy7FzFCxhMkepJscVJARoT8USR1PgNoSb1+upz+Q8POUb5IeljtM0+XY+gw
RvI4IKZrBYrLBJaK6TYm4fwu7r6p4xXXJUFLPDV5KLfpzoI3/qGbRtWKcHmoLS5X
Uk85NyqLBBkuGwLcyeokg4sG0YkEvQWDkFNvpcjIon++BfYHm77PMMytK0IpkGdp
lupS0V38MJNlW506NHG8TNcBPm3NBnjrk6qxfMEZGOWuk1+RUjCR3tNghEaaZ4gm
AbQEsRF23em0QtnfKqGImwvFC351ty0rXVDc0WhY3+J0DlRL9n5L9uu3ZQb1hE7z
c23AT8J2wQvgRKKerAn24alLE9WUgO92wioYmxBSVdMMgDgwaNCFCEDhOn/i2tNE
kMMlq3vAffPXoJJ7TWVP3MJm2Vtz5gUy0fsRXUaN1e+gFZ81QxPMseN0bRpa5P5r
diindpt+p1ob9JpZKgfpcXb1yDLUMF3u2RG4HxxB6ilcItKXQ22KzDPMk6Q3r2Gc
asNaJTcfoX3oDSCUMgxF0yBKwJlc3g1INZ613Nq2dRKuawW1y2LVgndeO7UcJazZ
NTIHmCzbm7kLnwzFHcVw81gGXomUppcxFn7oorq21dq9JRbRKj9mgoOrR5ZYDwhZ
c/rHXWhBUzeimGDa0BeUbojNYf2ykJNpMZCd5Xaw/9iOlSitW/hZ8gLqq/8Ul7fB
EHAPnLpW+nM1IyUastHaUmC4An5AIh4sPRrsS8rkqJttd02B+QsXE0Pw2tAbS2Up
is6Ffv3lRd4SHG6eJD+7R0MPiRwvw07ypEb5PFv8K6v68pVambbRvwLULilI2J6u
ICkHL58JOlMAzG7K4mecnT0y2LdW/eRmKyjIYE/PGKnSuKZT0YtBWX8wCKwI15L0
HzuhjxiABBtC5pLJZL0yTcMFu72JAAafv1QQuzYe8PGdMsCp4qw7Je762McjcHEs
1Ns7lhc64/23cal+xWsD8/QRkmfRurK8lgyXwRhHPWw1LX6k6F4cRmuLiYZGTN2m
dhhwHczgC08WXKqEr+siZQegBKLaHP/pLG17AVGn32hlAVCjPH8HsIGq61etSNMZ
dBtOQra8WNiKLZemiDsXVHG/OmSMvlmR/2foHQrqF/ouHRDkBoaDGIaa5Qw4N0Yk
aa+z3oKr05bLEJD7RoQO5lJhn+pI2tnjNUBSxtZxkIEi8Sii9CbLPF8mSyash8yD
tl7Vh39QlOpo4TdW1ajxRTe4IDyzAOTLvcaw+cv4P2liF8OEs2X/MveOYxKwXfUU
uk51e1pg0o3yJ5OJLu4CzqgTKmgNVV2MfoUDU++SEVl8uFhtxqsEGN/VfCe/IXJy
KieLFS1O+cJTN0T1R2Jhd25/EK6QUu217TctHlGzZVKJByPJ8S6rFqPetaQ/7edB
SShGObjEhAszi4LYUKdZmdgxzICdXvR/Xz6GmRJRzyHB6bxUhzZtIzka6uEUbvUd
tJkX2MHut8+/WitCVgb3OCE4Uf2FGRoe6lJ5A/zG0PfGfzuTl57bVX4zoGO36ic3
4YWcJ22+3Ggh1xWJhksofCMe5x/HNggnPFygT0tCJ331w+2OTkEYlcD6+jBRKQpE
m+kYkx7w/88Ljx2QS5/RQMgTev9ZcTVYVkBJPFtWmTZa8myBwVIRxcS7DNIf/+dY
+VMn7RLKLvs+/mO3tgxSb5G4eQdyhpUF7Da/f2IBBoy8xxmO/vA13iZwQLr1oIFc
VoyZh9z/T8DwBebxgzWyc16ki2mxucy6ZTREEH6MrPGu7V/u9v/F0do0M4EcIikd
unLHCJI2z64BEOrkIlzNwmK0+3Y0QsXfXp99n57ghG5XBGVZq2joGBGfbzdALnTy
Lr2aT8Qk172CgG0zOMgW3+4e2zj6eTrQN74zICB2BnW4ShnT7gr2HKK9ZlvKOQwO
IEDc+8BUZ6ZERXoKOhNLELsm8iRQ/Dpm7qO4cVwlsDHE47KvavUxSQIu1CP20Zea
LcTZhX/Q+b0g7NrgaN+NDDxY483AZHi4eXHUZHhrxBkM3iCsWw2zDEViB+Wm0WL9
0NecGPrqUfaJlH3crAP0wkLFdj7VN+2gnWSfL5vSxtUyGuiqxwO9DwaZOklqW62a
2WJMGbez+JlD0OE16AarqwMwMffNeFdwJxj81p/QQ2Fr66bmVE9/2QoXp3RNDGkO
qPvkbomGUoK7pXPTkwrZv+bNPiAAjGpEp/j4BYWfK6VDA5mAR8cpnIkfzoBehGWj
CeoULQ5pcFQYiQwUIx0JnWYXEkABGf6b0cb7Jqp5lzCPVxDbS4d6eiADbkPn+xWi
6AU0QRo/qVsYruB5IRBltauP0YuDbnN/xgzGf0BR9hMATZsKUChSrHPv2nzLkiEm
XR0DeaWsj6QpLJOpzZdnWuVTtdLof3L53yC/4/G3EBfkrL6XLellohZ0v/4RJmAy
ESfsXYfjFqb3J9Vdu805tdcECSE2Kj1lGOWtC5fLZ1DJdgSQe23RE/ZXol8vziKL
fr0BYeh/ScrwuaT6kK0VdUd2HTQLHFFXSZtvpuUkBD100UFhxgPxaJv28rwhm1Tx
xy45L9QUegfrYqcz4Ky1slPt/Dv0Q4AqDl9YnmRPfZMyTbMbEF1R5nUbRrZS4lC8
alIp9SgyySNCDXRlQZOaVJATf3YVnj7j4xuAL3G3fMG9kNtlL3PqR5OAvgXdeG/d
6sx1r1JTFPh8nf04obAECKBJJX+PL182TgWWH5Xrh5NB0g/ZrE09DmGR+RfL8yJA
4KQNTWxSr0vK+Bz9HCtenu/5clfCZPINwtY4R+KC4OYr7H8iUWm2f8ZKpBgDuNOR
fQRYX87BPcj4WrZAzcP2GUxPAWQjCtzlQRGcuYeXifL5VlucQFw9H+93lRuHTFDS
10EHrnRaAuQU0/Kn6lpL34TJs29mMmCNtgpQjbJo6mYtC4HfnNFL8oBe/BptRadv
CrPAPoKEvXEB1b1Bv+MKXWzmde2fWQA0N6qrG8IzcpXiW+kavoZ4d3RySxI03Xvc
Z65DyXjxEgFwKH1kWvEbT/bEqluzAyzho/St1xHmRSg7+KzaU+3JxPg9IOFGmTHA
BvZ8d79y4D4/xwntWfxkO/jjLIkEOKeEQMolY5XWCUo/ArbIovbYLI6AAH2os1xf
wgS7FYvaDUfVZQhgl8wECFO4VGa2QiiBMWv79HO4luxW7Fk7MZspAmbeCOKpW7a3
r5ZL38y2/x8ACjmWOxMNjTZu94ckSFkvU7i+xXPtFAFQ6caBCh2738CMR08x8iu1
4/HCzwE3vL8TRBY65pbuvldmLVjU7Wuv6FKIg2lFNGEusCNMEC19sZ69pkon6H3i
5QpZvGu32s1WgiexxB/e0KjbAjM8mkX3frhf2oUrGjPNMGTbeT1oex1E4E0yZbeN
CkbC4QPwFqF526uUfX07x6ZTqCGKEd8agAz4qrNoJ/wDVop/xZzlGTxAup6PTGMr
SjnbjKUjy7wt0dOQt11wmuz4WJQFjQ+OYuNJ/YTtfRGkb/d1lLirjaKOj2V1ngZe
qp+tJQhfIWWBsaZaqOvtdOIIVS5wNTVXakhPkcOYOLxyDEnvkdpVIDZVQWUV2vrr
5T3Z8ySl5fum7oLb356RXmV0CJf2COOQQgjaFRQSy+1QWrvnzymD//VReeTsUkfe
BvMGMLmO+0PFxvnKtrAlGbs7vWwt79QtWOymxckBQobOvnDqRIiPeCYIakhEY5rC
EqUXijttz4xKyORG32dg/Su6Gr5FHWcbvzgVMN8guWOJkUdaWsHVqqlvXiPrK6vL
Yl3aaPrMxwNm32+yxhbaUAW8jF2GNbGyK1Wd2X6HlNmcxwgSuTIyQFO7XbITyRl6
2Ws8U/qC7lORz0t7bF4tRtKSbuANmVYa7MFMIThqZtWKClz14Z6qTk51G9SDwe4E
IYtPZwK4V/G265NqCiZkgUHtYUzq+FEUFzPaFMRpZ79XujexXNokCw1ekSWvbIlR
7BtGMP/JN6WlPJa375rfGtEKu7Tstfhn8vcITCvmTe9M3t790R0TMZXHiOgyySCI
XIVKk7gZtNkZAV2A45cDtDIg85zAJB3K/WQsCxDUAzwkku9X6woIUa8pO+K/PdVv
8VgZk5q+6X3VCVoqsexvOcJ50h/BPmmso85/vBe+XHldKJohLiQSwH/iiesi8yM+
zUquRN7AyWnP1IEcZbBuv2slKu/p7Y6yj6npK4GR//gHLFXD5FeFQZIgV5e3EjMG
CJw6Pf8v7fNw4bZn1Qxdja+hiKzh6M8l8dVWqU/poipSAHHdMIgFYxWhUwYi2IsK
68hCBikxtUOEtEaYuVbLKo4axFhrDFAWlW06RAnooLaY6tQXjkyMRSmqIItg9jOe
SMNQHRdhoogn/xA6ed3G8Y3+UpWzxluBERhmf0FzyKeVqXnCK2LdN4wpgXTakmrZ
Sv2VY9LsaITvBG/mMRVjt6lntiAK9a8b1dtRt/+Ax/v58Qgc7nBxzdNSbufFgUdu
AexAFt1x+evgob21PIw6UsgWf1+nzv2jJs1ieUTPehtb4qDa4MoZ8CAkjbjtKcV3
x9L4aWDsNfKuY8o2UlzcEUPQjPSoq7RjtmDfSAhaHqUFv7ao5KguaMKS9m15r/Wb
N4pTSDY1PJySnO5eL9rVd6wJvuc/anOVZG8Ndxfzx9NZ0S24T9TDw/TdUCY7yc45
iNdUU187ENTyS54BAnpPjwvQ1mecwoPKnd48rCb8sIAjvh7eOCyazVYVkwH8Uu9k
AFqjiSh7Q/IUn36bgqKS07QS37ZmNuDZUNtKGXH9cVny9YbgXg+8MBczznyjo4ey
+rSvDfp6unkta9aEvHA1oMDr+EiRreBTIiznxifjn22kIkep2sksN2HzaSz8W2Sj
rZLX17Jvld4NiHNMH9INo5Rd+RtxpDm1KJxTc0L03V/sdEfMx2oSJklQoO25qvrw
bUgQZy5Uzf5SupLEYvcPy0CBHtleoAOekhwd2F4kwi/K4Y0CMRfOUW9CtcQXKoYV
n+FNfJcYuHR+whkuMfgdziRj9gl9BivTGPrpsHBCrhgZO9Cg3d3Zki5ECsD+beH9
zUdcxXKeNv4o/BOQCd+drVXgAZqQKwHTWTUaooRgTUYus2PQv2P4hfQXMjxOMtxc
IKuBLJnejW1SgTGTXIMQQes78CIAXL+1Ubod+0eQ4CV+32nGG+baxyGOs2NRZbyc
7tWQT818L7niiY7UsQcEZ50qVEPw22HHhC/xKTPksjiJ14e7pLyNtFIYUFeCI30P
8ERlISsuGP9UHYpnJV1OOdFYb2vl6TQxilB2Bl+AjXl1B4f/1ptrmolTkHYFAMob
AZFhqvmq9TDpNn9Lu0VlFHpOqTwpmSnFT0dQaB2clgketWC8OxbjxTszwOwfW5IR
OsLk7zHSTQB7JmFxnn1A6DEO1z/3ABj5CX5EaJd3YpVn50N7hrWUYpQJ4AMk3rxU
bPCX4vCGKDrH8H85MlgMVgPlKYhKwGDn22ZuvfckY2jyChwauXFUAiKHSbzIxo9+
CzQ+p2W5V0P0tGwXiCUC1xBvwKZCJIbacMbuqwO2nlurj/xV8OxX/uY1qTx3YHob
hMe5MfALv2GUoo9fcO5Vh/2ikXbW8LvlFNwnPHsEs4iWE/FNBlOXk8pF3zKSX18S
UyuAaOkYvwkgliK0MUNHbT7nWOcoZaD6BazkT6OjVT9gFjoslALPQRmOg3KBCZp8
qHzbcQVmaN3fhgJBRISdaphrIVlfMXAcQd7c3SlQWQri3MEZoXJcvej753YXUQr7
ZepRHUyMHt3LVnO1xVxRTHiGQmcpvxwuEuWaVbh9mzOpNf/8qvMkBxaYQK6S6Mj4
JnocwGNm9c3Ezx0UUv0wuOOX96S3ER9j2KZMm27a/vP7sQJMHVbHgFpbYIa+xREC
C359DU8QkGLUonWCLGxnXKsruNHh5Ie/ONEP65uqfgWoQXq8DaVgds2jIuK86j4z
wRoaX7MUkycOF5GPz/9YNthJoZ0PqbzXZziM+fmpPO98wrr2pmuY1CIQtu4M4aTG
3zK/THf16ytcNU1Rb57TTkMp9Mb6mTbV7iIJcS2aTkqHwOuTAaXsEApnu61GOgTI
iCiHYoZTq+1xhF2Wjofp9sJGxJkPaevP9NYBinWLcRzUhtNCrBH8RYdhbcLRABT7
zpY1tXoenN2pWCFDKsqSUDBEDVOQbAjvfuNg+P4JPUw4ntfKCafU4GI+Kyf75xn6
F8vrZtnNpmp93zF3BNV2l5EE0i0CFo5ByFCEu/bzkHC3gghuLb7F/yZM5eZbMD5x
sc0py7C5lSG8QtjTelRgFOP6bNrBg3XTW8IfxETJuoVwGTRsuOUDEN7l4bw8wWJA
oflblgA7iEku8mxw0jmkBbSEb3iPhsNW78McH/tolls8Ycii5oZbSIbOdnqtnmsH
1eozEoeT0NTQ1g/iLDtn8juRyPb3zIAFpGxaNDZMw9eH24010cNvLyIgsHyg7VLV
FEIhUoarljpOEDcn7ciqwl58QG5RDopKhiAD7o62QBP7NG1iBSURB8TLOpKbgd/c
`pragma protect end_protected



